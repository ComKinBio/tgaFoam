THERMO ALL
   300.000  1000.000  5000.000
AC3H4                   C   3H   4          G    300.00   3500.00 1800.00      1
 6.64430238e+00 1.14987825e-02-4.68099585e-06 9.62334222e-10-8.24360065e-14    2
 2.07131189e+04-1.35744541e+01 1.21562918e+00 2.35625008e-02-1.47340944e-05    3
 4.68570404e-09-5.99570704e-13 2.26674413e+04 1.58066578e+01                   4
ACETOL                  C   3H   6O   2     G    300.00   3500.00 1800.00      1
 9.43106557e+00 1.86879303e-02-7.29283976e-06 1.39932581e-09-1.08736168e-13    2
-4.87389994e+04-2.08360480e+01 1.41553145e+00 3.65002283e-02-2.21364215e-05    3
 6.89694866e-09-8.72294898e-13-4.58534071e+04 2.25456947e+01                   4
ALDEST                  C   6H  10O   3     G    300.00   3500.00 1800.00      1
 1.79608805e+01 3.27577303e-02-1.29904809e-05 2.50013680e-09-1.93431386e-13    2
-7.48983193e+04-5.99171462e+01 5.24137808e+00 6.10232913e-02-3.65451150e-05    3
 1.12240754e-08-1.40508952e-12-7.03192984e+04 8.92345431e+00                   4
ALDINS                  C  13H  20O   1     G    300.00   3500.00 1800.00      1
 8.44295858e+01 4.93170400e-02-2.86268350e-05 8.86979917e-09-1.00373619e-12    2
-8.94265291e+04-4.12065762e+02-1.18024916e+01 2.63166101e-01-2.06834386e-04    3
 7.48725957e-08-1.01707913e-11-5.47829813e+04 1.08762316e+02                   4
AR                      AR  1               G    300.00   3500.00 1490.00      1
 2.50000000e+00 7.40336223e-15-5.56967416e-18 1.73924876e-21-1.92673709e-25    2
-7.45375000e+02 4.36600000e+00 2.50000000e+00-4.07455160e-15 5.98527266e-18    3
-3.43074982e-21 6.74775716e-25-7.45375000e+02 4.36600000e+00                   4
BENZYNE                 C   6H   4          G    300.00   3500.00 1400.00      1
 1.09465819e+01 1.50373246e-02-5.27844959e-06 8.14607581e-10-4.49073366e-14    2
 5.03301418e+04-3.53782934e+01-3.73796173e+00 5.69931634e-02-5.02311341e-05    3
 2.22206478e-08-3.86741452e-12 5.44418140e+04 4.04070822e+01                   4
BIN1A                   C  20H  16          G    300.00   3500.00 1800.00      1
-3.24173600e+00 1.58222900e-01-9.46183500e-05 2.81843100e-08-3.56131000e-12    2
 2.17869900e+04 3.00825300e+01-3.24173600e+00 1.58222900e-01-9.46183500e-05    3
 2.81843100e-08-3.56131000e-12 2.17869900e+04 3.00825300e+01                   4
BIN1B                   C  20H  10          G    300.00   3500.00 1800.00      1
-5.70256700e+00 1.43432300e-01-8.80724700e-05 2.76799200e-08-3.52289900e-12    2
 2.77808900e+04 4.34481200e+01-5.70256700e+00 1.43432300e-01-8.80724700e-05    3
 2.76799200e-08-3.52289900e-12 2.77808900e+04 4.34481200e+01                   4
BIPHENYL                C  12H  10          G    300.00   3500.00 1450.00      1
 2.67692078e+01 2.81611415e-02-6.05667723e-06-3.69378426e-10 1.67249382e-13    2
 9.26692468e+03-1.21306413e+02-1.05625108e+01 1.31145193e-01-1.12591903e-04    3
 4.86123345e-08-8.27787353e-12 2.00931231e+04 7.26686556e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578334e+01 2.37623567e-02-8.52218599e-06 1.36123710e-09-7.97159891e-14    2
-5.90596972e+03-6.59480381e+01-8.70136947e+00 9.66875823e-02-8.77887356e-05    3
 3.96542562e-08-7.01685714e-12 1.03797027e+03 6.35339364e+01                   4
C                       C   1               G    300.00   3500.00  700.00      1
 2.48989675e+00 5.14965671e-05-7.37912415e-08 3.75721674e-11-4.86583734e-15    2
 8.54527782e+04 4.81783270e+00 2.55088394e+00-2.97001640e-04 6.72990632e-07    3
-6.73648664e-10 2.49141603e-13 8.54442400e+04 4.54535738e+00                   4
C10H10                  C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592698e+01 4.15934216e-02-1.83631832e-05 3.88491136e-09-3.27420808e-13    2
 4.39687821e+03-8.23923218e+01-1.14588964e+01 1.07633791e-01-7.33968243e-05    3
 2.42677414e-08-3.15836942e-12 1.50954180e+04 7.84485932e+01                   4
C10H6CH3                C  11H   9          G    300.00   3500.00 1800.00      1
 2.12659882e+01 3.44429430e-02-1.39605695e-05 2.72496148e-09-2.12674976e-13    2
 3.28507521e+04-9.11529083e+01-1.92673037e+00 8.59823175e-02-5.69100482e-05    3
 1.86321758e-08-2.42201030e-12 4.12001308e+04 3.43709226e+01                   4
C10H7                   C  10H   7          G    300.00   3500.00 1440.00      1
 1.86034915e+01 2.84557463e-02-7.51492092e-06 8.59843958e-11 1.31843536e-13    2
 3.89175328e+04-7.96671600e+01-8.11601745e+00 1.02676605e-01-8.48283149e-05    3
 3.58792224e-08-6.08226028e-12 4.66127513e+04 5.89821104e+01                   4
C10H7CH2                C  11H   9          G    300.00   3500.00 1460.00      1
 1.62958766e+01 4.54296741e-02-2.13529357e-05 4.77934912e-09-4.18010504e-13    2
 2.55100815e+04-6.47739136e+01-5.20583638e+00 1.04338477e-01-8.18756782e-05    3
 3.24153046e-08-5.15019466e-12 3.17885817e+04 4.70964540e+01                   4
C10H7CH3                C  11H  10          G    300.00   3500.00 1400.00      1
 1.59718633e+01 4.84656090e-02-2.27123224e-05 5.09437338e-09-4.47432797e-13    2
 5.32412011e+03-6.35417268e+01-7.85505905e+00 1.16542530e-01-9.56518805e-05    3
 3.98274963e-08-6.64977617e-12 1.19956584e+04 5.94264980e+01                   4
C10H7CHO                C  11H   8O   1     G    300.00   3500.00 1800.00      1
 2.76873866e+01 2.65153545e-02-9.85230690e-06 1.73492056e-09-1.21699947e-13    2
-1.08926269e+04-1.25645702e+02-1.80645208e+00 9.20572182e-02-6.44705267e-05    3
 2.19638908e-08-2.93127915e-12-2.74844971e+02 3.39811053e+01                   4
C10H7O                  C  10H   7O   1     G    300.00   3500.00 1800.00      1
 2.60845785e+01 2.24488808e-02-7.86244785e-06 1.25147148e-09-7.55452008e-14    2
 1.36168392e+03-1.17834769e+02-2.53985295e+00 8.60587284e-02-6.08706542e-05    3
 2.08841405e-08-2.80230479e-12 1.16664792e+04 3.70866255e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818224e+01 2.47079229e-02-8.75472975e-06 1.41213209e-09-8.61580367e-14    2
-1.58338687e+04-1.19314317e+02-3.09194614e+00 9.23929369e-02-6.74411581e-05    3
 2.40273261e-08-3.35424965e-12-5.70514482e+03 3.79602738e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248659e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987876e+01                   4
C11H12O4                C  11H  12O   4     G    300.00   3500.00 1280.00      1
 2.98957517e+01 4.73870505e-02-2.11603212e-05 4.60350399e-09-3.96349099e-13    2
-7.02119467e+04-1.21160681e+02-3.09348688e+00 1.50478421e-01-1.41970521e-04    3
 6.75254832e-08-1.26857982e-11-6.17667016e+04 4.61370519e+01                   4
C12H18                  C  12H  18          G    300.00   3500.00 1800.00      1
 8.44295858e+01 4.93170400e-02-2.86268350e-05 8.86979917e-09-1.00373619e-12    2
-8.94265291e+04-4.12065762e+02-1.18024916e+01 2.63166101e-01-2.06834386e-04    3
 7.48725957e-08-1.01707913e-11-5.47829813e+04 1.08762316e+02                   4
C12H22                  C  12H  22          G    300.00   3500.00 1760.00      1
 3.60687856e+01 4.93531801e-02-1.68932777e-05 2.64866878e-09-1.56934744e-13    2
-2.29291143e+04-1.58689972e+02-2.71855262e+00 1.37506222e-01-9.20237107e-05    3
 3.11071661e-08-4.19933494e-12-9.27597128e+03 5.03635315e+01                   4
C12H7                   C  12H   7          G    300.00   3500.00 1250.00      1
 1.23349807e+01 5.16907682e-02-2.72404819e-05 6.85858162e-09-6.72018930e-13    2
 5.30394981e+04-4.25244963e+01-8.02968441e+00 1.16857696e-01-1.05440796e-04    3
 4.85654157e-08-9.01338574e-12 5.81306643e+04 6.02674845e+01                   4
C12H8                   C  12H   8          G    300.00   3500.00 1430.00      1
 2.59652189e+01 2.42501190e-02-4.81412894e-06-4.21078741e-10 1.47447105e-13    2
 1.90778575e+04-1.18254954e+02-9.28199067e+00 1.22843712e-01-1.08233982e-04    3
 4.77933050e-08-8.28164096e-12 2.91585594e+04 6.43994840e+01                   4
C14H10                  C  14H  10          G    300.00   3500.00 1430.00      1
 3.13141255e+01 2.89528714e-02-5.57670990e-06-5.89662906e-10 1.88202945e-13    2
 1.06460191e+04-1.48101025e+02-1.21905872e+01 1.50644375e-01-1.33225141e-04    3
 5.89200950e-08-1.02156009e-11 2.30883669e+04 7.73445897e+01                   4
C14H9                   C  14H   9          G    300.00   3500.00 1430.00      1
 3.13141255e+01 2.89528714e-02-5.57670990e-06-5.89662906e-10 1.88202945e-13    2
 4.06560892e+04-1.48101025e+02-1.21905872e+01 1.50644375e-01-1.33225141e-04    3
 5.89200950e-08-1.02156009e-11 5.30984370e+04 7.73445897e+01                   4
C16H10                  C  16H  10          G    300.00   3500.00 1430.00      1
 3.55205969e+01 2.97059226e-02-5.18577408e-06-7.74976601e-10 2.05764301e-13    2
 1.13998034e+04-1.72584653e+02-1.43149515e+01 1.69106058e-01-1.51409692e-04    3
 6.73946823e-08-1.17120082e-11 2.56527702e+04 8.56679628e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933977e+01 6.96117135e-02-3.71054121e-05 9.43826014e-09-9.32515880e-13    2
 4.61008358e+04-6.54256237e+01-1.33382684e+01 1.64875153e-01-1.52343443e-04    3
 7.13941909e-08-1.34236310e-11 5.34246890e+04 8.34001920e+01                   4
C2-OOQOOH               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323243e+01 1.62358927e-02-6.84260319e-06 1.39267431e-09-1.12911127e-13    2
-1.87641105e+04-2.90906767e+01 5.81911522e+00 3.09319129e-02-1.90892866e-05    3
 5.92848300e-09-7.42884555e-13-1.63833552e+04 6.70139036e+00                   4
C2-OQOOH                C   2H   4O   3     G    300.00   3500.00 1800.00      1
 1.06961666e+01 1.25934013e-02-5.32391821e-06 1.08565058e-09-8.80671200e-14    2
-3.42000230e+04-2.43964294e+01 5.53941294e+00 2.40528540e-02-1.48734621e-05    3
 4.62251869e-09-5.79298801e-13-3.23435917e+04 3.51299738e+00                   4
C2-QOOH                 C   2H   5O   2     G    300.00   3500.00 1270.00      1
 7.85685775e+00 1.67911217e-02-7.79621720e-06 1.73782470e-09-1.51982948e-13    2
 7.20248835e+02-1.06887184e+01 8.24295798e-01 3.89409231e-02-3.39574000e-05    3
 1.54707291e-08-2.85531058e-12 2.50651957e+03 2.49202290e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1770.00      1
 2.62706056e+00 5.61439161e-03-2.33738366e-06 4.29433761e-10-2.92352464e-14    2
 6.73836200e+04 9.73315238e+00 4.71151838e+00 9.03752455e-04 1.65468342e-06    3
-1.07416966e-09 1.83138118e-13 6.66457220e+04-1.51333448e+00                   4
C2H2                    C   2H   2          G    300.00   3500.00  970.00      1
 4.61193612e+00 5.01498204e-03-1.65253694e-06 2.49922532e-10-1.30568636e-14    2
 2.56043843e+04-3.75517096e+00 1.83812159e+00 1.64533925e-02-1.93408005e-05    3
 1.24068047e-08-3.14627391e-12 2.61425043e+04 9.54239252e+00                   4
C2H2O2                  C   2H   2O   2     G    300.00   3500.00 1700.00      1
 9.83116579e+00 4.87360532e-03-1.69443300e-06 2.65361078e-10-1.54439841e-14    2
-2.96273239e+04-2.66407027e+01 1.89947966e+00 2.35363962e-02-1.81616014e-05    3
 6.72307419e-09-9.65107677e-13-2.69305506e+04 1.58338747e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00  700.00      1
 7.05094230e-01 1.53761148e-02-8.91788178e-06 2.51340905e-09-2.70561650e-13    2
 3.36189510e+04 1.96531878e+01 2.74606708e+00 3.71341276e-03 1.60736225e-05    3
-2.12880236e-08 8.22995002e-12 3.33332148e+04 1.05346375e+01                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1340.00      1
 6.70517760e+00 1.61222451e-02-7.57298869e-06 1.70307233e-09-1.49924851e-13    2
-1.33618589e+04-9.88613663e+00 3.40917666e-01 3.51200360e-02-2.88391725e-05    3
 1.22832633e-08-2.12384107e-12-1.16562372e+04 2.26803642e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1800.00      1
 4.49333672e+00 1.00335105e-02-3.62601388e-06 5.97613541e-10-3.65481279e-14    2
 3.93220822e+03-3.35192020e+00 2.66161697e-01 1.94272328e-02-1.14541158e-05    3
 3.49691054e-09-4.39228267e-13 5.45399123e+03 1.95264329e+01                   4
C2H4CHO                 C   3H   5O   1     G    300.00   3500.00  760.00      1
 2.15579434e+00 2.57531407e-02-1.33069384e-05 3.28122872e-09-3.12828174e-13    2
-7.31459492e+02 1.94816815e+01 3.58641615e+00 1.82235522e-02 1.55409151e-06    3
-9.75476244e-09 3.97532681e-12-9.48914007e+02 1.29723736e+01                   4
C2H4O                   C   2H   4O   1     G    300.00   3500.00 1440.00      1
 4.77217531e+00 1.29608883e-02-4.19608017e-06 3.32859470e-10 2.97428516e-14    2
-8.91054882e+03-2.99568268e+00-1.76683146e+00 3.11247960e-02-2.31168173e-05    3
 9.09246001e-09-1.49102113e-12-7.02731487e+03 3.09356489e+01                   4
C2H4O2                  C   2H   4O   2     G    300.00   3500.00  770.00      1
 3.40614010e+00 2.02613044e-02-1.03463461e-05 2.53497107e-09-2.40436915e-13    2
-3.88060356e+04 1.20569218e+01 4.64403525e+00 1.38306802e-02 2.18084389e-06    3
-8.31108086e-09 3.28100852e-12-3.89966715e+04 6.40833543e+00                   4
C2H4OH                  C   2H   5O   1     G    300.00   3500.00 1800.00      1
 6.43071837e+00 1.30529032e-02-5.04234033e-06 9.42421880e-10-7.06192378e-14    2
-6.84254175e+03-6.40643970e+00 1.19058412e+00 2.46976460e-02-1.47462926e-05    3
 4.53647829e-09-5.69793739e-13-4.95609342e+03 2.19542600e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00  700.00      1
-1.10489358e+00 2.43511913e-02-1.39613152e-05 3.89870297e-09-4.17285120e-13    2
 1.35030749e+04 3.00146907e+01 4.99501831e+00-1.05054480e-02 6.07314834e-05    3
-6.72372957e-08 2.49884287e-11 1.26490872e+04 2.76182763e+00                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1140.00      1
-3.19796156e+00 4.17401347e-02-2.22156952e-05 5.37596466e-09-4.95601240e-13    2
-2.31457657e+04 4.43385409e+01 4.65967589e+00 1.41694770e-02 1.40614860e-05    3
-1.58387612e-08 4.15675092e-12-2.49373071e+04 5.40040975e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1380.00      1
 4.82959470e+00 1.77552121e-02-6.21112100e-06 6.58265206e-10 1.60136692e-14    2
-3.08658494e+04 5.43180378e-01 2.48921589e-01 3.10325255e-02-2.06429833e-05    3
 7.63017938e-09-1.24701426e-12-2.96015836e+04 2.41176395e+01                   4
C2H5OO                  C   2H   5O   2     G    300.00   3500.00 1260.00      1
 4.82335647e+00 2.06819188e-02-9.67611879e-06 2.17589519e-09-1.91914821e-13    2
-4.75156327e+03 3.93765088e+00 1.82119985e+00 3.02125747e-02-2.10221378e-05    3
 8.17907984e-09-1.38302289e-12-3.99501980e+03 1.91151548e+01                   4
C2H5OOH                 C   2H   6O   2     G    300.00   3500.00 1590.00      1
 1.15652199e+01 1.02216474e-02-1.86630047e-06-2.55692055e-10 7.26211298e-14    2
-2.47328137e+04-3.42112965e+01 1.46294225e+00 3.56361824e-02-2.58422768e-05    3
 9.79712822e-09-1.50801099e-12-2.15202894e+04 1.92111233e+01                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.39373503e+00 1.52684734e-02-5.82725051e-06 1.10377088e-09-8.60486537e-14    2
-1.27269866e+04-3.21997495e+00-2.74461309e-01 2.56422430e-02-1.44720586e-05    3
 4.30555164e-09-5.30740425e-13-1.10464360e+04 2.20452775e+01                   4
C3-OQOOH                C   3H   6O   3     G    300.00   3500.00 1350.00      1
 1.12132537e+01 2.34709018e-02-1.13098317e-05 2.59008079e-09-2.30885268e-13    2
-3.91289882e+04-2.66260028e+01 8.46220448e-01 5.41880374e-02-4.54399824e-05    3
 1.94444762e-08-3.35206960e-12-3.63298893e+04 2.65001343e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00  700.00      1
 6.27665898e+00 5.58433105e-03-2.45857473e-06 5.41223006e-10-4.83608105e-14    2
 6.31055207e+04-4.75111128e+00 4.26055345e+00 1.71049341e-02-2.71455812e-05    3
 2.40526578e-08-8.44530180e-12 6.33877755e+04 4.25633816e+00                   4
C3H3                    C   3H   3          G    300.00   3500.00 1720.00      1
 1.09930471e+01 7.79714852e-04 1.73957383e-06-7.95864951e-10 9.69732207e-14    2
 3.74627231e+04-3.40822737e+01 3.56039712e+00 1.80649474e-02-1.33347569e-05    3
 5.04689889e-09-7.52265710e-13 4.00195547e+04 5.80687271e+00                   4
C3H4O2                  C   3H   4O   2     G    300.00   3500.00 1240.00      1
 1.02920429e+01 1.38871300e-02-6.12561993e-06 1.30548845e-09-1.09965765e-13    2
-3.57026988e+04-2.69350036e+01 1.17378045e-01 4.67086294e-02-4.58290467e-05    3
 2.26514168e-08-4.41358036e-12-3.31793820e+04 2.43405589e+01                   4
C3H4O3                  C   3H   4O   3     G    300.00   3500.00 1710.00      1
 1.37242810e+01 1.08811110e-02-3.70124855e-06 5.78901440e-10-3.43205818e-14    2
-5.77802807e+04-3.99570073e+01 2.17563103e+00 3.78954970e-02-2.73980784e-05    3
 9.81743159e-09-1.38498288e-12-5.38306424e+04 2.19543274e+01                   4
C3H5CHO                 C   4H   6O   1     G    300.00   3500.00 1610.00      1
 9.36564259e+00 1.99394689e-02-8.24714277e-06 1.63840913e-09-1.29181894e-13    2
-1.44293663e+04-2.07054000e+01 2.40474771e-01 4.26106933e-02-2.93694015e-05    3
 1.03846860e-08-1.48729943e-12-1.14910622e+04 2.76639767e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00  820.00      1
 2.45863176e+00 2.66446458e-02-1.24879759e-05 2.92198798e-09-2.71872686e-13    2
-1.72239991e+04 1.83830345e+01 4.24999286e+00 1.79062989e-02 3.49680492e-06    3
-1.00737688e-08 3.69024828e-12-1.75177823e+04 1.00962500e+01                   4
C3H5OO                  C   3H   5O   2     G    300.00   3500.00 1800.00      1
 7.69230110e+00 2.05361077e-02-9.61589847e-06 2.15332094e-09-1.88909485e-13    2
 6.21484234e+03-1.04053755e+01 2.96424215e+00 3.10429054e-02-1.83715632e-05    3
 5.39615972e-09-6.39303761e-13 7.91694356e+03 1.51838658e+01                   4
C3H5OOH                 C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.21377197e+01 1.68585481e-02-6.94275126e-06 1.36958900e-09-1.07427460e-13    2
-1.25265904e+04-3.57194708e+01 2.24651097e+00 3.88390118e-02-2.52598044e-05    3
 8.15368275e-09-1.04966270e-12-8.96575529e+03 1.78138141e+01                   4
C3H6                    C   3H   6          G    300.00   3500.00 1800.00      1
 9.21549195e+00 1.10096151e-02-2.72165887e-06 1.69301120e-10 1.25058839e-14    2
-2.15028535e+03-2.75773224e+01-2.61886761e-01 3.20704567e-02-2.02723602e-05    3
 6.66956086e-09-8.90307969e-13 1.26157099e+03 2.37162283e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1720.00      1
 6.42754902e+00 2.00818525e-02-6.55464685e-06 4.84306793e-10 5.68893699e-14    2
-1.48035725e+04-9.71995026e+00-9.99780843e-02 3.52621481e-02-1.97932767e-05    3
 5.61555868e-09-6.88932126e-13-1.25581031e+04 2.53116313e+01                   4
C3H6O2                  C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.08721654e+01 1.63593216e-02-6.08637842e-06 1.10130850e-09-8.02911326e-14    2
-4.55272952e+04-2.70748520e+01 2.66105929e+00 3.46062241e-02-2.12921305e-05    3
 6.73306853e-09-8.62480026e-13-4.25712970e+04 1.73653673e+01                   4
C3H7CHO                 C   4H   8O   1     G    300.00   3500.00  700.00      1
-9.77279434e-01 5.24983747e-02-3.09762338e-05 8.32680251e-09-8.38156520e-13    2
-2.70767712e+04 3.27194912e+01 3.71554492e+00 2.56822356e-02 2.64869216e-05    3
-4.64000121e-08 1.87071344e-11-2.77337666e+04 1.17531393e+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   3500.00 1670.00      1
 1.20273024e+01 2.23669330e-02-9.25510611e-06 1.83134653e-09-1.43510571e-13    2
-2.87878078e+04-3.43698022e+01 1.14029559e+00 4.84435961e-02-3.26772586e-05    3
 1.11815072e-08-1.54323522e-12-2.51515476e+04 2.37368269e+01                   4
C3H8                    C   3H   8          G    300.00   3500.00 1800.00      1
 1.08596364e+01 1.35766563e-02-3.19926248e-06 1.41615801e-10 2.35898562e-14    2
-1.80884704e+04-3.69486914e+01-1.25512725e+00 4.04983533e-02-2.56340099e-05    3
 8.45078153e-09-1.13046094e-12-1.37271555e+04 2.86189366e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00 1050.00      1
 8.50275797e+00 6.97445022e-03-2.53297106e-06 4.33287765e-10-2.93611469e-14    2
 5.31727553e+04-2.08807943e+01 2.90907865e+00 2.82837048e-02-3.29747633e-05    3
 1.97614098e-08-4.63129497e-12 5.43474279e+04 6.37839155e+00                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208969e+01 1.53590365e-03 1.80568199e-06-9.30237202e-10 1.18077197e-13    2
 6.01811751e+04-4.25791500e+01 2.34662667e+00 2.83894138e-02-2.35278181e-05    3
 9.69177542e-09-1.55205057e-12 6.35755930e+04 1.38680560e+01                   4
C4H3O                   C   4H   3O   1     G    300.00   3500.00 1240.00      1
 8.44125905e+00 1.62911136e-02-8.34126436e-06 2.01436766e-09-1.87394603e-13    2
 1.94535776e+04-2.27855078e+01-5.90872253e+00 6.25813767e-02-6.43375505e-05    3
 3.21198978e-08-6.25705794e-12 2.30123730e+04 4.95317026e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1190.00      1
 6.36293592e+00 1.66610000e-02-7.54220850e-06 1.59521425e-09-1.28415834e-13    2
 3.13137240e+04-8.19255288e+00 4.03184847e-01 3.66937767e-02-3.27936077e-05    3
 1.57416564e-08-3.10035746e-12 3.27321448e+04 2.15965194e+01                   4
C4H4O                   C   4H   4O   1     G    300.00   3500.00 1250.00      1
 8.37486466e+00 1.95634451e-02-9.90167121e-06 2.37694382e-09-2.20517698e-13    2
-9.41817580e+03-2.52053384e+01-7.59507781e+00 7.06672610e-02-7.12262503e-05    3
 3.50833860e-08-6.76180613e-12-5.42569018e+03 5.54039922e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794385e-03 4.88814513e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742307e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H6                    C   4H   6          G    300.00   3500.00 1550.00      1
 9.55395345e+00 1.51364811e-02-4.78509457e-06 6.14955374e-10-2.23809938e-14    2
 8.63284693e+03-2.77966685e+01-1.04533857e+00 4.24894928e-02-3.12557510e-05    3
 1.20001840e-08-1.85870818e-12 1.19186275e+04 2.79839806e+01                   4
C4H6O2                  C   4H   6O   2     G    300.00   3500.00 1800.00      1
 7.01919581e+00 2.89919962e-02-1.39811163e-05 3.22750474e-09-2.90888810e-13    2
-4.36055710e+04-7.47846940e+00 9.15158242e-01 4.25565241e-02-2.52848896e-05    3
 7.41408744e-09-8.72358628e-13-4.14081175e+04 2.55578553e+01                   4
C4H7OH                  C   4H   8O   1     G    300.00   3500.00 1460.00      1
 1.00981665e+01 2.15734935e-02-6.74008418e-06 9.16825971e-10-4.16200161e-14    2
-2.37290909e+04-2.45741592e+01-2.55531336e-01 4.99397889e-02-3.58835384e-05    3
 1.42243393e-08-2.32030381e-12-2.07058111e+04 2.92946643e+01                   4
C4H8O                   C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.12815996e+01 2.48463701e-02-1.13234700e-05 2.47069946e-09-2.12413507e-13    2
-2.03756688e+04-3.84267373e+01-2.94845122e+00 5.64687053e-02-3.76754160e-05    3
 1.22306795e-08-1.56796629e-12-1.52528505e+04 3.85892666e+01                   4
C4H9CHO                 C   5H  10O   1     G    300.00   3500.00  760.00      1
-1.78433179e+00 6.31204386e-02-3.60836198e-05 9.48321920e-09-9.39522544e-13    2
-2.97113508e+04 3.92478712e+01 5.53299014e+00 2.46082180e-02 3.99273421e-05    3
-5.71930632e-08 2.09934651e-11-3.08235837e+04 5.95416540e+00                   4
C4H9OOH                 C   4H  10O   2     G    300.00   3500.00 1780.00      1
 1.73966948e+01 2.30088698e-02-8.34646932e-06 1.39883190e-09-9.01677555e-14    2
-3.38614042e+04-6.23628946e+01 1.12895120e+00 5.95655969e-02-3.91527000e-05    3
 1.29367460e-08-1.71066131e-12-2.80700874e+04 2.54997628e+01                   4
C5EN-OO                 C   5H   9O   2     G    300.00   3500.00 1280.00      1
 1.00840321e+01 3.69913036e-02-1.74216180e-05 3.93130749e-09-3.47257402e-13    2
-8.98415155e+02-1.96513637e+01 4.09897281e-01 6.72229749e-02-5.28493577e-05    3
 2.23832553e-08-3.95115346e-12 1.57816336e+03 2.94089022e+01                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   3500.00 1160.00      1
 1.36699765e+01 4.21231935e-02-2.15503712e-05 5.21806336e-09-4.87293014e-13    2
-1.42354804e+04-3.35883364e+01 5.24578583e-01 8.74521518e-02-8.01654035e-05    3
 3.89048635e-08-7.74737926e-12-1.11857480e+04 3.17816498e+01                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   3500.00 1580.00      1
 1.69833146e+01 2.73095032e-02-1.19226853e-05 2.48166925e-09-2.03420392e-13    2
-3.51234520e+04-5.58041780e+01 1.44561329e+00 6.66454559e-02-4.92669442e-05    3
 1.82387405e-08-2.69662788e-12-3.02135384e+04 2.62635800e+01                   4
C5EN-QOOH               C   5H   9O   2     G    300.00   3500.00 1420.00      1
 1.28791275e+01 3.32930454e-02-1.55378924e-05 3.46674396e-09-3.02869803e-13    2
 3.23011716e+03-3.38507184e+01 1.34404411e+00 6.57862381e-02-4.98616876e-05    3
 1.95812018e-08-3.13992224e-12 6.50608085e+03 2.58442475e+01                   4
C5H4O2                  C   5H   4O   2     G    300.00   3500.00 1430.00      1
 1.05158962e+01 2.23224229e-02-1.09267096e-05 2.56683236e-09-2.34844997e-13    2
-2.33303219e+04-2.94000374e+01-1.81996644e+00 5.68283325e-02-4.71217197e-05    3
 1.94409629e-08-3.18486782e-12-1.98022652e+04 3.45255921e+01                   4
C5H5O                   C   5H   5O   1     G    300.00   3500.00 1450.00      1
 1.05801390e+01 2.13128784e-02-9.63052935e-06 2.09384798e-09-1.79321204e-13    2
 1.62543411e+04-3.26154734e+01-4.01979397e+00 6.15885556e-02-5.12950230e-05    3
 2.12499370e-08-3.48209517e-12 2.04883217e+04 4.32455666e+01                   4
C5H7                    C   5H   7          G    300.00   3500.00 1430.00      1
 7.72404525e+00 2.56072196e-02-8.76350316e-06 8.66193959e-10 3.30416650e-14    2
 2.30808142e+04-1.69352935e+01 2.31765047e-01 4.65646468e-02-3.07468184e-05    3
 1.11148258e-08-1.75867718e-12 2.52236063e+04 2.18904247e+01                   4
C5H8                    C   5H   8          G    300.00   3500.00 1430.00      1
 8.95829159e+00 2.51033002e-02-8.43679234e-06 8.19905621e-10 3.11426511e-14    2
 4.67953300e+03-2.40439628e+01 1.19183502e+00 4.68276543e-02-3.12245763e-05    3
 1.14435811e-08-1.82614328e-12 6.90073958e+03 1.62025638e+01                   4
C5H8O                   C   5H   8O   1     G    300.00   3500.00 1330.00      1
 6.70800688e+00 3.65243775e-02-1.77765821e-05 4.15639148e-09-3.79163309e-13    2
-5.52771782e+03-9.67918417e+00-5.12640161e+00 7.21165834e-02-5.79181678e-05    3
 2.42774871e-08-4.16132413e-12-2.37976516e+03 5.07899199e+01                   4
C5H8O4                  C   5H   8O   4     G    300.00   3500.00 1230.00      1
 1.19601536e+01 3.99450843e-02-1.95947373e-05 4.60940117e-09-4.22302290e-13    2
-8.26385858e+04-2.91875208e+01-6.95683231e+00 1.01463738e-01-9.46174851e-05    3
 4.52721371e-08-8.68708602e-12-7.79850073e+04 6.59920851e+01                   4
C5H9CHO                 C   6H  10O   1     G    300.00   3500.00 1800.00      1
 1.08416239e+01 4.20296686e-02-2.00742994e-05 4.57927363e-09-4.08519043e-13    2
-3.59631714e+04-3.80017802e+01-6.51363638e+00 8.05969136e-02-5.22136702e-05    3
 1.64827443e-08-2.06177886e-12-2.97152777e+04 5.59285088e+01                   4
C6H10O5                 C   6H  10O   5     G    300.00   3500.00 1220.00      1
 1.54889718e+01 4.96354387e-02-2.45944509e-05 5.82332585e-09-5.35665863e-13    2
-1.09180509e+05-4.81819837e+01-7.95116461e+00 1.26488345e-01-1.19085729e-04    3
 5.74579042e-08-1.11165221e-11-1.03461116e+05 6.95642163e+01                   4
C6H2                    C   6H   2          G    300.00   3500.00 1100.00      1
 1.20007067e+01 9.35747205e-03-3.45039279e-06 5.96931921e-10-4.08067421e-14    2
 8.10797696e+04-3.61630610e+01 4.40206371e+00 3.69889013e-02-4.11296144e-05    3
 2.34328238e-08-5.23078218e-12 8.27514710e+04 1.22022725e+00                   4
C6H3                    C   6H   3          G    300.00   3500.00 1320.00      1
 1.19194523e+01 1.16137832e-02-4.19264523e-06 6.84693072e-10-4.17887568e-14    2
 8.26280760e+04-3.29876543e+01 4.46601450e+00 3.41999583e-02-2.98587533e-05    3
 1.36473739e-08-2.49684195e-12 8.45957836e+04 5.04018537e+00                   4
C6H4                    C   6H   4          G    300.00   3500.00 1360.00      1
 1.74447675e+01 6.21306708e-03-9.80963858e-07 8.00594635e-11-2.88320770e-15    2
 5.49568894e+04-6.59208082e+01-1.17305610e+00 6.09713718e-02-6.13761529e-05    3
 2.96855443e-08-5.44506791e-12 6.00209374e+04 2.96241244e+01                   4
C6H4C2H                 C   8H   5          G    300.00   3500.00 1490.00      1
 3.21415686e+01-1.98168404e-02 2.64282529e-05-1.09843473e-08 1.50630597e-12    2
 5.44964091e+04-1.47026437e+02-4.78252619e+00 7.93082463e-02-7.33621030e-05    3
 3.36645815e-08-5.98512503e-12 6.54997893e+04 4.58354239e+01                   4
C6H4CH3                 C   7H   7          G    300.00   3500.00 1450.00      1
 1.23344954e+01 2.38147082e-02-7.01721971e-06 3.58622104e-10 7.92842393e-14    2
 2.97091697e+04-3.94240761e+01-4.14387803e+00 6.92722902e-02-5.40423045e-05    3
 2.19793508e-08-3.64842760e-12 3.44878980e+04 4.61973136e+01                   4
C6H4O2                  C   6H   4O   2     G    300.00   3500.00 1410.00      1
 1.74929577e+01 1.29021286e-02-2.02976642e-06-3.72417846e-10 8.59745727e-14    2
-2.22100459e+04-6.49015838e+01-5.23446578e+00 7.73770890e-02-7.06201498e-05    3
 3.20580235e-08-5.66410367e-12-1.58009124e+04 5.25540058e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1690.00      1
 2.37494889e+01-3.74826288e-03 7.22829016e-06-2.69927706e-09 3.10032681e-13    2
 2.93571719e+04-1.07010346e+02-4.30972117e+00 6.26640688e-02-5.17175663e-05    3
 2.05535263e-08-3.12973113e-12 3.88411849e+04 4.30825907e+01                   4
C6H5C2H                 C   8H   6          G    300.00   3500.00 1330.00      1
 1.36301627e+01 2.67826138e-02-1.18276978e-05 2.56807250e-09-2.21616638e-13    2
 3.04381476e+04-4.83434869e+01-3.73085925e+00 7.89962135e-02-7.07152163e-05    3
 3.20856256e-08-5.77002888e-12 3.50561794e+04 4.03644060e+01                   4
C6H5C2H2                C   8H   7          G    300.00   3500.00 1690.00      1
 1.77155600e+01 2.19043174e-02-8.07391246e-06 1.39474201e-09-9.41524347e-14    2
 3.81394494e+04-7.01114193e+01-2.50848763e+00 6.97718858e-02-5.05599199e-05    3
 1.81545083e-08-2.57340780e-12 4.49751775e+04 3.80700548e+01                   4
C6H5C2H3                C   8H   8          G    300.00   3500.00 1420.00      1
 1.57612121e+01 2.51344730e-02-7.08348959e-06 3.12355848e-10 8.22985790e-14    2
 1.01346894e+04-5.95859946e+01-4.61890423e+00 8.25432514e-02-6.77265654e-05    3
 2.87832834e-08-4.93018867e-12 1.59226425e+04 4.58827137e+01                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   3500.00 1440.00      1
 2.29999925e+01 5.23551496e-02-1.62023052e-05 1.06346924e-09 1.48747565e-13    2
 3.20131872e+03-9.18704227e+01-1.05589612e+01 1.45574466e-01-1.13305759e-04    3
 4.60187721e-08-7.65599251e-12 1.28662974e+04 8.22691715e+01                   4
C6H5C2H5                C   8H  10          G    300.00   3500.00 1440.00      1
 1.53992430e+01 3.11284429e-02-9.32920034e-06 5.29654938e-10 9.71609974e-14    2
-4.32725762e+03-5.77491740e+01-6.11786341e+00 9.08981829e-02-7.15893461e-05    3
 2.93537965e-08-4.90703025e-12 1.86966902e+03 5.39044909e+01                   4
C6H5CH2C6H5             C  13H  12          G    300.00   3500.00 1440.00      1
 2.36600260e+01 4.20961068e-02-1.18756749e-05 4.02369975e-10 1.68531444e-13    2
 4.50897730e+03-9.76688099e+01-1.18613481e+01 1.40766591e-01-1.14657429e-04    3
 4.79865153e-08-8.09260490e-12 1.47391331e+04 8.66539117e+01                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799879e-06 4.38368241e-10 8.64078959e-14    2
-1.87828963e+04-3.81332333e+01-6.02884975e+00 7.77532977e-02-6.10481840e-05    3
 2.48568442e-08-4.12367417e-12-1.33857950e+04 5.85676633e+01                   4
C6H5CHO                 C   7H   6O   1     G    300.00   3500.00 1770.00      1
 2.73588480e+01 2.45725463e-03 5.41130341e-06-2.58531717e-09 3.21649872e-13    2
-1.76429542e+04-1.23608292e+02-6.55705980e+00 7.91033740e-02-5.95430351e-05    3
 2.18795937e-08-3.13384602e-12-5.63672287e+03 5.93816475e+01                   4
C6H5O                   C   6H   5O   1     G    300.00   3500.00 1320.00      1
 1.34428169e+01 1.79658729e-02-6.67332779e-06 1.12237517e-09-7.10809502e-14    2
 4.07683820e+02-4.72500520e+01-4.80707078e+00 7.32685627e-02-6.95172935e-05    3
 3.28617518e-08-6.08232652e-12 5.22565416e+03 4.58618544e+01                   4
C6H5OCH3                C   7H   8O   1     G    300.00   3500.00 1380.00      1
 1.25085136e+01 3.49906122e-02-1.63096082e-05 3.64836832e-09-3.19988393e-13    2
-1.52038795e+04-4.20406499e+01-5.29461551e+00 8.65938851e-02-7.24001222e-05    3
 3.07452350e-08-5.22884105e-12-1.02902159e+04 4.95832512e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1330.00      1
 1.39867712e+01 2.02277643e-02-7.36599500e-06 1.21196288e-09-7.46105018e-14    2
-1.80542263e+04-5.08485811e+01-5.47325435e+00 7.87541571e-02-7.33732049e-05    3
 3.42982836e-08-6.29384372e-12-1.28778595e+04 4.85843830e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1550.00      1
 1.57365829e+01 1.24444139e-02-2.08242468e-06-1.90555168e-10 5.60938650e-14    2
 2.37538837e+03-6.60380946e+01-6.33361145e+00 6.93997541e-02-5.72004958e-05    3
 2.35161421e-08-3.76756698e-12 9.21714860e+03 5.01102066e+01                   4
C6H6O3                  C   6H   6O   3     G    300.00   3500.00 1770.00      1
 1.98638073e+01 1.79335016e-02-5.95408859e-06 8.93593939e-10-4.95459880e-14    2
-4.95264845e+04-7.44496694e+01 7.10718582e-01 6.12173180e-02-4.26352889e-05    3
 1.47094886e-08-2.00094354e-12-4.27462910e+04 2.88889342e+01                   4
C6H8O4                  C   6H   8O   4     G    300.00   3500.00 1300.00      1
 1.58073709e+01 3.77998882e-02-1.77241312e-05 3.97560136e-09-3.49009860e-13    2
-7.78788467e+04-5.15128322e+01-4.55493836e+00 1.00453147e-01-9.00163533e-05    3
 4.10485358e-08-7.47842033e-12-7.25846463e+04 5.20658817e+01                   4
C7DIONE                 C   7H  12O   2     G    300.00   3500.00  700.00      1
-7.55853587e-01 8.24536116e-02-4.58824665e-05 1.18274999e-08-1.15807940e-12    2
-3.67546790e+04 2.64722477e+01 3.52180397e+00 5.80098541e-02 6.49701379e-06    3
-3.80577194e-08 1.66580704e-11-3.73535510e+04 7.36075600e+00                   4
C7H15COCHO              C   9H  16O   2     G    300.00   3500.00 1780.00      1
 3.02050983e+01 3.84107591e-02-1.30454122e-05 2.02881682e-09-1.19348346e-13    2
-6.67956450e+04-1.25747051e+02 3.59041588e-01 1.05480549e-01-6.95648985e-05    3
 2.31971638e-08-3.09243078e-12-5.61704488e+04 3.54525548e+01                   4
C7H7                    C   7H   7          G    300.00   3500.00 1450.00      1
 1.55564029e+01 1.97467971e-02-4.90102499e-06-1.06746050e-11 9.16513058e-14    2
 1.67098727e+04-6.15086686e+01-4.40172355e+00 7.48036976e-02-6.18564392e-05    3
 2.61757227e-08-4.42324479e-12 2.24977294e+04 4.21934668e+01                   4
C7H8                    C   7H   8          G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799879e-06 4.38368241e-10 8.64078959e-14    2
-5.64471283e+02-4.45247833e+01-6.02884975e+00 7.77532977e-02-6.10481840e-05    3
 2.48568442e-08-4.12367417e-12 4.83263000e+03 5.21761133e+01                   4
C7KETONE                C   7H  14O   1     G    300.00   3500.00 1800.00      1
 1.82994273e+01 4.14393597e-02-1.71834162e-05 3.42714287e-09-2.72037363e-13    2
-4.27848802e+04-6.59785823e+01-2.29236271e-01 8.26141675e-02-5.14957561e-05    3
 1.61354169e-08-2.03707542e-12-3.61145614e+04 3.43024100e+01                   4
C8H10O3                 C   8H  10O   3     G    300.00   3500.00 1280.00      1
 2.98957517e+01 4.73870505e-02-2.11603212e-05 4.60350399e-09-3.96349099e-13    2
-7.02119467e+04-1.21160681e+02-3.09348688e+00 1.50478421e-01-1.41970521e-04    3
 6.75254832e-08-1.26857982e-11-6.17667016e+04 4.61370519e+01                   4
C8H2                    C   8H   2          G    300.00   3500.00 1060.00      1
 1.62719352e+01 9.99874492e-03-2.93037080e-06 2.89537341e-10 2.52405898e-16    2
 1.07885460e+05-5.89733614e+01 1.87361722e-01 7.06952484e-02-8.88216494e-05    3
 5.43092094e-08-1.27402363e-11 1.11295389e+05 1.95626382e+01                   4
C8H9                    C   8H   9          G    300.00   3500.00 1570.00      1
 2.45973914e+01 1.20503967e-02 5.66754133e-07-1.10955314e-09 1.57308310e-13    2
 1.65948730e+04-1.06442126e+02-5.12604623e+00 8.77789001e-02-7.17853192e-05    3
 2.96131956e-08-4.73484913e-12 2.59280324e+04 5.03637968e+01                   4
C9H10O2                 C   9H  10O   2     G    300.00   3500.00 1620.00      1
 2.64048781e+01 2.84903123e-02-1.03289369e-05 1.78607618e-09-1.22280426e-13    2
-3.71439509e+04-1.10770565e+02-2.04331024e+00 9.87327525e-02-7.53682334e-05    3
 2.85512188e-08-4.25270367e-12-2.79267379e+04 4.01996488e+01                   4
CH                      C   1H   1          G    300.00   3500.00 1720.00      1
 1.56762354e+00 3.35441204e-03-1.29971595e-06 2.40500907e-10-1.78141164e-14    2
 7.11686733e+04 1.27712404e+01 3.85901271e+00-1.97439999e-03 3.34750385e-06    3
-1.56074708e-09 2.43995183e-13 7.03804355e+04 4.73936215e-01                   4
CH2                     C   1H   2          G    300.00   3500.00  900.00      1
 3.24505871e+00 2.75395076e-03-7.68471343e-07 8.23040037e-11-1.89900250e-15    2
 4.54794580e+04 4.28187007e+00 3.99717917e+00-5.88806826e-04 4.80279129e-06    3
-4.04455721e-09 1.14445133e-12 4.53440763e+04 7.32567433e-01                   4
CH2C3H5                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45916998e+00 1.93968541e-02-5.99075606e-06 3.82147973e-10 5.73994806e-14    2
 1.98988324e+04-1.80212793e+01-3.29329051e-01 4.23733221e-02-2.85167051e-05    3
 1.01973763e-08-1.54639600e-12 2.25881131e+04 2.81156134e+01                   4
CH2CCH3                 C   3H   5          G    300.00   3500.00 1800.00      1
 1.00124373e+01 7.55815802e-03-1.17096962e-06-2.01794819e-10 4.72987983e-14    2
 2.78641947e+04-2.75169832e+01 6.10512020e-01 2.84513252e-02-1.85819423e-05    3
 6.24671358e-09-8.48327368e-13 3.12488878e+04 2.33681976e+01                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   3500.00 1590.00      1
 1.05858550e+01 1.29956017e-02-4.76361255e-06 7.49449815e-10-3.96847802e-14    2
 3.10513348e+03-2.93262371e+01 1.05972039e+00 3.69607201e-02-2.73722149e-05    3
 1.02289476e-08-1.53017186e-12 6.13444428e+03 2.10494483e+01                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.17572858e+01 2.41574264e-02-9.72976868e-06 1.89143875e-09-1.46945289e-13    2
-1.45672160e+04-3.14377946e+01 8.93764133e-01 4.82985857e-02-2.98474014e-05    3
 9.34241382e-09-1.18180294e-12-1.06563482e+04 2.73578508e+01                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   3500.00 1800.00      1
 9.49770379e+00 1.77061096e-02-6.68456978e-06 1.20981994e-09-8.73179586e-14    2
-1.07976200e+04-2.07829255e+01 1.04629052e+00 3.64870279e-02-2.23353351e-05    3
 7.00639969e-09-8.92398479e-13-7.75511123e+03 2.49578861e+01                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097165e-06 1.27900113e-09-8.37238502e-14    2
-1.74897435e+04-4.46134901e+01 9.11733056e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH2CHCH2                C   3H   5          G    300.00   3500.00 1800.00      1
 1.31270112e+01 3.37812631e-03 1.30787951e-06-8.72502093e-10 1.13779857e-13    2
 1.38569110e+04-4.71985703e+01 1.45788193e-01 3.22252886e-02-2.27314224e-05    3
 8.03094306e-09-1.12280975e-12 1.85301513e+04 2.30585168e+01                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   3500.00 1780.00      1
 1.38129918e+01 2.02819032e-02-7.03372780e-06 1.12439860e-09-6.86002896e-14    2
-1.64045579e+04-4.42517079e+01 2.32452600e-01 5.07999690e-02-3.27511989e-05    3
 1.07564103e-08-1.42141092e-12-1.15698860e+04 2.90972641e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1030.00      1
 3.66502520e+00 1.44768244e-02-7.23266377e-06 1.70580456e-09-1.56345856e-13    2
-3.68579193e+01 5.92341850e+00 2.15742069e-01 2.78720987e-02-2.67403448e-05    3
 1.43321353e-08-3.22098924e-12 6.73694406e+02 2.26661724e+01                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   3500.00 1380.00      1
 6.32694430e+00 2.38762490e-02-1.07376178e-05 2.33737032e-09-2.01069469e-13    2
-1.14217376e+04-3.95690500e+00 6.40756935e-01 4.03579515e-02-2.86525118e-05    3
 1.09919085e-08-1.76892059e-12-9.85234986e+03 2.53070892e+01                   4
CH2CHOOHCHO             C   3H   5O   3     G    300.00   3500.00 1300.00      1
 1.09154411e+01 2.11069264e-02-1.04347901e-05 2.43633157e-09-2.20224944e-13    2
-1.35446352e+04-2.42468452e+01 1.81101363e+00 4.91205495e-02-4.27582013e-05    3
 1.90124399e-08-3.40793808e-12-1.11774841e+04 2.20654311e+01                   4
CH2CN                   C   2H   2N   1     G    300.00   3500.00  980.00      1
 4.41880974e+00 9.83430327e-03-4.98991807e-06 1.22319871e-09-1.17396557e-13    2
 2.92390343e+04 2.02769260e+00 2.71162977e+00 1.68023848e-02-1.56553489e-05    3
 8.47859386e-09-1.96826267e-12 2.95736416e+04 1.02293594e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1410.00      1
 6.03578795e+00 5.81722422e-03-1.93206512e-06 2.83140054e-10-1.50051612e-14    2
-8.58422380e+03-7.64505060e+00 2.49197065e+00 1.58706066e-02-1.26271528e-05    3
 5.33991909e-09-9.11597189e-13-7.58486732e+03 1.06694385e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  930.00      1
 1.06639253e+00 1.06960337e-02-5.54447373e-06 1.36053696e-09-1.28442554e-13    2
-1.46324373e+04 1.74071779e+01 3.13463322e+00 1.80037482e-03 8.80336316e-06    3
-8.92465077e-09 2.63639286e-12-1.50171301e+04 7.57920580e+00                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1590.00      1
 7.61004151e+00 1.40239019e-03 1.05265418e-06-5.61972284e-10 7.11209072e-14    2
-5.04985629e+03-1.55757586e+01 1.95857131e+00 1.56199253e-02-1.23601148e-05    3
 5.06183022e-09-8.13124769e-13-3.25268877e+03 1.43100973e+01                   4
CH2OOCH2CHO             C   3H   5O   3     G    300.00   3500.00 1800.00      1
 1.06998539e+01 2.42793089e-02-1.34097218e-05 3.42673974e-09-3.32159552e-13    2
-2.14126656e+04-2.48508794e+01 2.93009251e+00 4.15454454e-02-2.77981689e-05    3
 8.75579421e-09-1.07230601e-12-1.86155515e+04 1.72006902e+01                   4
CH2OOCHOOHCHO           C   3H   5O   5     G    300.00   3500.00 1800.00      1
 2.14549192e+01 1.08256409e-02-3.75393277e-06 5.88014009e-10-3.47282962e-14    2
-3.59900210e+04-7.93559883e+01 5.41191662e+00 4.64767576e-02-3.34631967e-05    3
 1.15914451e-08-1.56298261e-12-3.02145401e+04 7.47208818e+00                   4
CH2OOHCHCHO             C   3H   5O   3     G    300.00   3500.00  700.00      1
 1.84816700e+00 3.99042619e-02-2.38947704e-05 6.48850081e-09-6.57628290e-13    2
-1.48991977e+04 2.15340498e+01 5.44326670e+00 1.93608350e-02 2.01268587e-05    3
-3.54368602e-08 1.43157149e-11-1.54025117e+04 5.47205385e+00                   4
CH2OOHCHOOCHO           C   3H   5O   5     G    300.00   3500.00 1800.00      1
 2.14549192e+01 1.08256409e-02-3.75393277e-06 5.88014009e-10-3.47282962e-14    2
-3.59900210e+04-7.93559883e+01 5.41191662e+00 4.64767576e-02-3.34631967e-05    3
 1.15914451e-08-1.56298261e-12-3.02145401e+04 7.47208818e+00                   4
CH2S                    C   1H   2          G    300.00   3500.00  900.00      1
 2.57518275e+00 4.11179659e-03-1.68232435e-06 3.44404948e-10-2.93085968e-14    2
 5.01958500e+04 6.99914504e+00 4.62572654e+00-5.00173140e-03 1.35068890e-05    3
-1.09068642e-08 3.09604394e-12 4.98267521e+04-2.67749711e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1270.00      1
 2.57723974e+00 6.62601164e-03-2.54906392e-06 4.67320141e-10-3.34867663e-14    2
 1.65488693e+04 6.94195966e+00 3.53327401e+00 3.61488008e-03 1.00739068e-06    3
-1.39958516e-09 3.34014277e-13 1.63060366e+04 2.10113860e+00                   4
CH3C10H6O               C  11H   9O   1     G    300.00   3500.00 1800.00      1
 2.60936624e+01 3.24954978e-02-1.30480618e-05 2.52260906e-09-1.95492396e-13    2
-2.87396993e+03-1.14905139e+02-1.85059487e+00 9.45938472e-02-6.47966864e-05    3
 2.16887663e-08-2.85745868e-12 7.18596268e+03 3.63350107e+01                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   3500.00 1800.00      1
 2.91191869e+01 2.86451308e-02-9.80098219e-06 1.51374083e-09-8.72237944e-14    2
-2.13626711e+04-1.32660114e+02-1.76841814e+00 9.72842531e-02-6.70002508e-05    3
 2.26986551e-08-3.02957300e-12-1.02431333e+04 3.45100483e+01                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   3500.00  700.00      1
 2.02076663e+00 4.09903683e-02-2.06486866e-05 5.00507647e-09-4.71523451e-13    2
-1.40718373e+04 2.15880986e+01 3.53447938e+00 3.23405812e-02-2.11342851e-06    3
-1.26475503e-08 5.83298611e-12-1.42837571e+04 1.48252130e+01                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.16093380e+01 2.56981798e-02-1.09676558e-05 2.25993093e-09-1.85313976e-13    2
-1.31948148e+04-3.43573902e+01 5.90549372e-02 5.13654755e-02-3.23570689e-05    3
 1.01819358e-08-1.28559243e-12-9.03671291e+03 2.81551514e+01                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.30151659e+01 2.21750012e-02-8.49156594e-06 1.54860371e-09-1.12013678e-13    2
-1.79081220e+04-4.01994427e+01 1.75489331e+00 4.71978292e-02-2.93439226e-05    3
 9.27169878e-09-1.18466577e-12-1.38544238e+04 2.07435017e+01                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 9.07749584e+00 1.96975457e-02-8.18089073e-06 1.64328968e-09-1.31786153e-13    2
-9.31061125e+03-2.21687275e+01 2.91958855e-01 3.92209612e-02-2.44504037e-05    3
 7.66903521e-09-9.68695255e-13-6.14781793e+03 2.53804314e+01                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.15124775e+01 2.41072597e-02-9.86401997e-06 1.98674692e-09-1.62119892e-13    2
-1.58991633e+04-3.03580006e+01 1.53457350e-01 4.93495266e-02-3.08992425e-05    3
 9.77757006e-09-1.24417866e-12-1.18099160e+04 3.11193861e+01                   4
CH3CH2CHOCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.30434362e+01 2.38164771e-02-9.82552432e-06 1.93897534e-09-1.51918988e-13    2
-1.58538336e+04-4.35088383e+01 4.17731726e-02 5.27090615e-02-3.39026780e-05    3
 1.08564397e-08-1.39045570e-12-1.11732349e+04 2.68588742e+01                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   3500.00 1620.00      1
 8.28181025e+00 2.00744959e-02-8.21041648e-06 1.62349331e-09-1.27917758e-13    2
-1.30492834e+04-1.56179098e+01 1.73835403e+00 3.62311779e-02-2.31703072e-05    3
 7.77982697e-09-1.07796925e-12-1.09292035e+04 1.91072184e+01                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097165e-06 1.27900113e-09-8.37238502e-14    2
-1.74897435e+04-4.46134901e+01 9.11733056e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   3500.00 1430.00      1
 8.72382272e+00 3.04342830e-02-1.39185549e-05 3.06043861e-09-2.64689231e-13    2
-1.80661273e+04-1.71435098e+01 1.27395834e+00 5.12730645e-02-3.57774166e-05    3
 1.32510501e-08-2.04626467e-12-1.59354661e+04 2.14624055e+01                   4
CH3CH3-C5H6             C   7H  12          G    300.00   3500.00 1310.00      1
 1.53755546e+01 3.27318283e-02-1.05955708e-05 1.52102630e-09-7.69415914e-14    2
-6.19682930e+03-5.37226046e+01-1.29247813e+00 8.36265847e-02-6.88720094e-05    3
 3.11782470e-08-5.73671653e-12-1.82980473e+03 3.11918393e+01                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.15124775e+01 2.41072597e-02-9.86401997e-06 1.98674692e-09-1.62119892e-13    2
-1.58991633e+04-3.03580006e+01 1.53457350e-01 4.93495266e-02-3.08992425e-05    3
 9.77757006e-09-1.24417866e-12-1.18099160e+04 3.11193861e+01                   4
CH3CHCH2OCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.38488385e+01 2.14834842e-02-8.03028843e-06 1.42167056e-09-9.95437051e-14    2
-1.51249440e+04-4.82209549e+01-4.69026374e-01 5.33009618e-02-3.45448531e-05    3
 1.12418797e-08-1.46346164e-12-9.97051265e+03 2.92703168e+01                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 7.64501934e+00 2.06996931e-02-8.77824684e-06 1.84245353e-09-1.55992331e-13    2
-1.15050426e+04-1.08131884e+01 5.39035202e-01 3.64907690e-02-2.19374767e-05    3
 6.71624238e-09-8.32907449e-13-8.94688828e+03 2.76458802e+01                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   3500.00 1450.00      1
 8.91411879e+00 2.94184843e-02-1.30488503e-05 2.81020956e-09-2.39749810e-13    2
-1.71145335e+04-1.85255698e+01 6.16106328e-01 5.23095531e-02-3.67292664e-05    3
 1.36977572e-08-2.11691319e-12-1.47081099e+04 2.45907827e+01                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.11524016e+01 2.52912378e-02-1.05179486e-05 2.12392650e-09-1.71553011e-13    2
-1.78095410e+04-2.94209720e+01 6.76902371e-01 4.85701251e-02-2.99170213e-05    3
 9.30876825e-09-1.16944770e-12-1.40383613e+04 2.72746153e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.27018126e+00 1.06201871e-02-3.82264672e-06 6.56340789e-10-4.60549581e-14    2
-2.29794782e+04-8.60119259e+00 9.91751377e-01 2.23500313e-02-1.35975169e-05    3
 4.27666307e-09-5.48877497e-13-2.10792434e+04 1.99667711e+01                   4
CH3CHOH                 C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.00303702e+00 2.30237358e-02-1.19372743e-05 2.98274467e-09-2.88183748e-13    2
-6.17751011e+03 2.39401608e+01 1.83915526e+00 1.82459173e-02-1.69909177e-06    3
-6.76790535e-09 3.19419126e-12-6.29456667e+03 2.02045961e+01                   4
CH3CHOOCHO              C   3H   5O   3     G    300.00   3500.00 1800.00      1
 1.58771657e+01 1.28699615e-02-5.29703385e-06 1.04001953e-09-8.12487153e-14    2
-2.38887629e+04-5.44666587e+01 3.38301196e+00 4.06347476e-02-2.84343556e-05    3
 9.60939795e-09-1.27144016e-12-1.93908676e+04 1.31543077e+01                   4
CH3CN                   C   2H   3N   1     G    300.00   3500.00  700.00      1
 2.02660925e+00 1.64402545e-02-8.54290907e-06 2.13740318e-09-2.08581596e-13    2
 8.61823027e+03 1.31030643e+01 2.36621609e+00 1.44996440e-02-4.38445795e-06    3
-1.82302645e-09 1.20585756e-12 8.57068531e+03 1.15857868e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 5.59449005e+00 8.95063669e-03-3.42706569e-06 6.39554414e-10-4.91680987e-14    2
-5.31931220e+03-3.46466160e+00 1.83189171e+00 1.73119663e-02-1.03948404e-05    3
 3.22021171e-09-4.07592723e-13-3.96477680e+03 1.68993055e+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469381e+01 2.48483421e-03 1.65900438e-06-8.55133987e-10 9.82287242e-14    2
-2.73756816e+04-4.36816972e+01 2.64892548e+00 2.83894083e-02-2.04187576e-05    3
 7.50765465e-09-1.08966739e-12-2.33635811e+04 1.77505788e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1760.00      1
 1.54960865e+01 1.58758106e-03 2.24425901e-06-9.74237206e-10 1.03773065e-13    2
-4.69655432e+04-5.18401164e+01 3.62388957e+00 2.85698467e-02-2.07519902e-05    3
 7.73646324e-09-1.13354234e-12-4.27865299e+04 1.21478877e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 9.24187097e+00 1.34946785e-02-5.23722666e-06 9.72748882e-10-7.19834442e-14    2
-8.04571079e+03-2.24258259e+01 1.82620860e+00 2.99739283e-02-1.89699348e-05    3
 6.05893707e-09-7.78398470e-13-5.37607233e+03 1.77092859e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00  700.00      1
 8.22157368e-01 3.18964631e-02-1.68324056e-05 4.20706053e-09-4.04124926e-13    2
-2.74737271e+04 2.17873546e+01 1.03654018e+00 3.06714184e-02-1.42073099e-05    3
 1.70696939e-09 4.88764769e-13-2.75037407e+04 2.08295464e+01                   4
CH3COHCH3               C   3H   7O   1     G    300.00   3500.00 1270.00      1
 6.71652579e+00 2.35306498e-02-1.06144747e-05 2.31761627e-09-1.99886320e-13    2
-1.44175086e+04-7.90476332e+00 1.21649821e+00 4.08535713e-02-3.10746182e-05    3
 1.30578491e-08-2.31410538e-12-1.30205016e+04 1.99442900e+01                   4
CH3COOH                 C   2H   4O   2     G    300.00   3500.00 1410.00      1
 7.83491620e+00 1.12357063e-02-3.13558070e-06 1.59502818e-10 3.01357560e-14    2
-5.57414981e+04-1.53809923e+01 3.13168541e-01 3.25739975e-02-2.58358905e-05    3
 1.08925098e-08-1.87287967e-12-5.36203653e+04 2.34914872e+01                   4
CH3NO                   C   1H   3O   1N   1G    300.00   3500.00  860.00      1
 1.73828229e+00 1.65479495e-02-8.69271695e-06 2.17002760e-09-2.08463444e-13    2
 8.36473513e+03 1.74966005e+01 2.23451684e+00 1.42398818e-02-4.66701756e-06    3
-9.50669597e-10 6.98715974e-13 8.27938279e+03 1.51773992e+01                   4
CH3NO2                  C   1H   3O   2N   1G    300.00   3500.00 1620.00      1
 5.94771391e+00 1.22319078e-02-4.98716389e-06 9.73177561e-10-7.54873508e-14    2
-1.14691242e+04-2.73415041e+00-2.05952276e-01 2.74261453e-02-1.90559023e-05    3
 6.76278185e-09-9.68944802e-13-9.47533640e+03 2.99224212e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00  700.00      1
 6.88420582e-01 1.44971301e-02-7.59068052e-06 1.92522389e-09-1.90011116e-13    2
 1.18330404e+03 1.95838279e+01 2.13962537e+00 6.20453130e-03 1.01791740e-05    3
-1.49984471e-08 5.85415708e-12 9.80135371e+02 1.31002120e+01                   4
CH3OCH2                 C   2H   5O   1     G    300.00   3500.00  750.00      1
 2.76373432e+00 2.09427776e-02-1.03906311e-05 2.45853855e-09-2.25935821e-13    2
-6.59718889e+02 1.23154396e+01 2.98724171e+00 1.97507382e-02-8.00655224e-06    3
 3.39357381e-10 4.80457902e-13-6.93244997e+02 1.13014447e+01                   4
CH3OCH3                 C   2H   6O   1     G    300.00   3500.00  700.00      1
 8.15389478e-01 2.72675400e-02-1.40181429e-05 3.43685384e-09-3.25542356e-13    2
-2.31745898e+04 1.99239256e+01 1.74097325e+00 2.19784899e-02-2.68446400e-06    3
-7.35712603e-09 3.52945045e-12-2.33041715e+04 1.57886515e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 2.14769740e+00 2.46740524e-02-1.35238094e-05 3.44782067e-09-3.34980467e-13    2
-4.40372636e+04 1.69024645e+01 3.51192337e+00 1.68784755e-02 3.18099831e-06    3
-1.24615200e-08 5.34692693e-12-4.42282552e+04 1.08074480e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849390e-09-3.11411020e-13    2
-2.07085510e+04 1.59117693e+01 4.66126893e+00 9.68655554e-03 1.14715528e-05    3
-1.83003965e-08 7.03409939e-12-2.10131064e+04 6.50453092e+00                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00  700.00      1
 9.34193000e-01 1.60266556e-02-8.00101466e-06 1.97129714e-09-1.91599484e-13    2
-2.50979789e+04 1.91008457e+01 2.88895785e+00 4.85657077e-03 1.59348814e-05    3
-2.08247943e-08 7.94986176e-12-2.53716460e+04 1.03674509e+01                   4
CH3ONO                  C   1H   3O   2N   1G    300.00   3500.00 1800.00      1
 8.58034518e+00 8.90954082e-03-3.35922089e-06 6.18588139e-10-4.68096982e-14    2
-1.15569624e+04-1.97194056e+01 1.99249583e+00 2.35492060e-02-1.55589419e-05    3
 5.13700333e-09-6.74367363e-13-9.18533663e+03 1.59354094e+01                   4
CH3ONO2                 C   1H   3O   3N   1G    300.00   3500.00 1800.00      1
 1.07457798e+01 1.03362024e-02-4.39539782e-06 8.95959797e-10-7.26862027e-14    2
-1.81031090e+04-3.08875015e+01 1.35155390e+00 3.12122600e-02-2.17921125e-05    3
 7.33918744e-09-9.67578931e-13-1.47211877e+04 1.99560088e+01                   4
CH3OO                   C   1H   3O   2     G    300.00   3500.00 1300.00      1
 3.46521970e+00 1.23938518e-02-5.59614682e-06 1.22616716e-09-1.06238815e-13    2
 6.86982281e+02 1.04298931e+01 4.30117244e+00 9.82168948e-03-2.62826727e-06    3
-2.95822349e-10 1.86451475e-13 4.69634569e+02 6.17758023e+00                   4
CH3OOH                  C   1H   4O   2     G    300.00   3500.00 1800.00      1
 5.50146514e+00 1.13975421e-02-3.82130848e-06 4.38704910e-10-2.90617476e-15    2
-1.79784234e+04-4.65581411e-01 5.93430876e+00 1.04356674e-02-3.01974623e-06    3
 1.41830001e-10 3.83264515e-14-1.81342471e+04-2.80822136e+00                   4
CH4                     C   1H   4          G    300.00   3500.00 1070.00      1
-2.82321416e-01 1.42739336e-02-6.77628877e-06 1.55380951e-09-1.39473841e-13    2
-9.36383584e+03 2.03507024e+01 2.85765313e+00 2.53571100e-03 9.67916346e-06    3
-8.69880870e-09 2.25599770e-12-1.00357904e+04 4.98969392e+00                   4
CHCHCH3                 C   3H   5          G    300.00   3500.00 1800.00      1
 1.00124373e+01 7.55815802e-03-1.17096962e-06-2.01794819e-10 4.72987983e-14    2
 2.78641947e+04-2.75169832e+01 6.10512020e-01 2.84513252e-02-1.85819423e-05    3
 6.24671358e-09-8.48327368e-13 3.12488878e+04 2.33681976e+01                   4
CN                      C   1N   1          G    300.00   3500.00  810.00      1
 2.73859606e+00 2.23580966e-03-1.33797023e-06 4.34996429e-10-5.05222621e-14    2
 5.14568835e+04 8.20480076e+00 4.08532688e+00-4.41471288e-03 1.09778123e-05    3
-9.70145006e-09 3.07801060e-12 5.12387131e+04 1.99138758e+00                   4
CO                      C   1O   1          G    300.00   3500.00 1000.00      1
 2.68595014e+00 2.12486373e-03-1.04548608e-06 2.45538864e-10-2.22550981e-14    2
-1.41423615e+04 7.96579426e+00 3.81890943e+00-2.40697343e-03 5.75226966e-06    3
-4.28629830e-09 1.11070419e-12-1.43689533e+04 2.49992060e+00                   4
CO2                     C   1O   2          G    300.00   3500.00 1620.00      1
 5.07830985e+00 2.05366041e-03-5.94311265e-07 5.38675131e-11 1.66346855e-15    2
-4.92442103e+04-4.47815290e+00 2.44892797e+00 8.54596135e-03-6.60570102e-06    3
 2.52769046e-09-3.80099332e-13-4.83922906e+04 9.47557732e+00                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673687e+01 3.34155283e-02-1.38949871e-05 2.56768166e-09-1.71519559e-13    2
-2.17187243e+04-3.95715124e+01-4.41843936e+00 8.43645604e-02-7.22335735e-05    3
 3.22565297e-08-5.83733025e-12-1.73470426e+04 4.54334869e+01                   4
CSOLID                  C   1               S    300.00   3500.00 1470.00      1
 1.73007911e+00 1.24133836e-03-3.99676695e-07 5.50148663e-11-1.79078883e-15    2
-8.17038240e+02-1.00735633e+01-8.82758554e-01 8.35110072e-03-7.65453624e-06    3
 3.34520060e-09-5.61346186e-13-4.88639663e+01 3.53849619e+00                   4
CYC5H4O                 C   5H   4O   1     G    300.00   3500.00 1260.00      1
 6.34459579e+00 2.39841575e-02-8.32755388e-06 8.47127653e-10 2.86249484e-14    2
 3.08659308e+03-9.73181554e+00-5.14379339e+00 6.04552342e-02-5.17455024e-05    3
 2.38195872e-08-4.52940274e-12 5.98166715e+03 4.83481227e+01                   4
CYC5H5                  C   5H   5          G    300.00   3500.00  700.00      1
 4.01652575e+00 2.68451891e-02-1.26423018e-05 2.78092332e-09-2.35299436e-13    2
 2.91110159e+04 1.44025794e+00-2.58737408e+00 6.45817595e-02-9.35063814e-05    3
 7.97943325e-08-2.77400884e-11 3.00355619e+04 3.09448116e+01                   4
CYC5H6                  C   5H   6          G    300.00   3500.00 1020.00      1
 1.70141558e+00 3.79065957e-02-2.19495256e-05 6.12706526e-09-6.63672518e-13    2
 1.38484401e+04 1.22453451e+01-6.32922867e+00 6.93993183e-02-6.82623529e-05    3
 3.63968870e-08-8.08274648e-12 1.54866915e+04 5.11475893e+01                   4
CYC5H8                  C   5H   8          G    300.00   3500.00 1460.00      1
 8.43099915e+00 2.71082714e-02-1.07932862e-05 1.95387666e-09-1.31111174e-13    2
-1.09862538e+03-2.37608447e+01-6.56863980e+00 6.82031726e-02-5.30140751e-05    3
 2.12327757e-08-3.43229252e-12 3.28126920e+03 5.42801525e+01                   4
CYC6-OO                 C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.87814621e+01 3.54361927e-02-1.49718784e-05 3.04328287e-09-2.46478319e-13    2
-1.95252830e+04-7.87240875e+01-6.50623568e+00 9.16310766e-02-6.18009483e-05    3
 2.03873828e-08-2.65538109e-12-1.04217118e+04 5.81382079e+01                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283791e-14    2
-3.55499047e+04-1.29752781e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.56593329e+01                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283791e-14    2
-3.55499047e+04-1.29752781e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.56593329e+01                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283791e-14    2
-3.55499047e+04-1.30447295e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.49648189e+01                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.17655243e+01 3.67451404e-02-1.42717448e-05 2.74140449e-09-2.13135508e-13    2
-3.59903393e+04-5.10812501e+01-1.06696444e+01 9.82113560e-02-7.74219664e-05    3
 3.15771221e-08-5.15075839e-12-2.94392700e+04 6.56457555e+01                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415883e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.91587814e+01-8.02402159e+00 8.95009509e-02-6.86853396e-05    3
 2.77298318e-08-4.50893790e-12-3.06512867e+04 5.29538877e+01                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415883e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.98532958e+01-8.02402159e+00 8.95009509e-02-6.86853396e-05    3
 2.77298318e-08-4.50893790e-12-3.06512867e+04 5.22593733e+01                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.91384147e+01 3.64873063e-02-1.63612962e-05 3.53264562e-09-3.02111689e-13    2
-1.43294351e+04-7.86383640e+01-4.87015408e+00 8.98396814e-02-6.08216088e-05    3
 1.99994281e-08-2.58916481e-12-5.68635037e+03 5.13010187e+01                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300723e+01 3.28719793e-02-1.40160778e-05 2.89193638e-09-2.38539838e-13    2
-1.52994543e+04-8.89349636e+01-7.04914219e+00 9.50480115e-02-6.58294380e-05    3
 2.20820698e-08-2.90383614e-12-5.22693704e+03 6.24943819e+01                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300723e+01 3.28719793e-02-1.40160778e-05 2.89193638e-09-2.38539838e-13    2
-1.52994543e+04-8.89349636e+01-7.04914219e+00 9.50480115e-02-6.58294380e-05    3
 2.20820698e-08-2.90383614e-12-5.22693704e+03 6.24943819e+01                   4
CYC6H10                 C   6H  10          G    300.00   3500.00 1800.00      1
 1.51624858e+01 2.76360017e-02-1.05259858e-05 1.89586361e-09-1.35054773e-13    2
-9.29985245e+03-6.25064559e+01-6.01517655e+00 7.46974737e-02-4.97438791e-05    3
 1.64210093e-08-2.15243611e-12-1.67589399e+03 5.21114707e+01                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.29323176e+01 2.20056554e-02-7.35242348e-06 1.07816406e-09-5.64635915e-14    2
-2.79806200e+04-1.10525204e+02-1.05629257e+01 9.64395294e-02-6.93806518e-05    3
 2.40515820e-08-3.24721608e-12-1.59223324e+04 7.07580407e+01                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.18028612e+01 2.41377428e-02-8.73118284e-06 1.46035609e-09-9.51866870e-14    2
-2.87387454e+04-1.06217525e+02-1.25990095e+01 1.00586344e-01-7.24383509e-05    3
 2.50556035e-08-3.37230438e-12-1.63540719e+04 7.99725758e+01                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.14079592e+01 2.50825461e-02-9.38039634e-06 1.64525432e-09-1.14247640e-13    2
-3.89741817e+04-1.05728233e+02-1.45960517e+01 1.05091459e-01-7.60544907e-05    3
 2.63393633e-08-3.54398500e-12-2.60127378e+04 8.91329846e+01                   4
CYC6H10-ONE             C   6H  10O   1     G    300.00   3500.00 1800.00      1
 1.15965428e+01 4.02887933e-02-1.86685839e-05 4.15568433e-09-3.64030709e-13    2
-3.62221493e+04-4.27468434e+01-6.46490379e+00 8.04253413e-02-5.21157073e-05    3
 1.65435078e-08-2.08456175e-12-2.97200285e+04 5.50054734e+01                   4
CYC6H11                 C   6H  11          G    300.00   3500.00 1800.00      1
 1.12879190e+01 3.94798364e-02-1.80474738e-05 3.97976998e-09-3.47933573e-13    2
 4.69934406e+02-4.15743644e+01-9.20200373e+00 8.50129981e-02-5.59917752e-05    3
 1.80332150e-08-2.29980093e-12 7.84630661e+03 6.93213721e+01                   4
CYC6H12                 C   6H  12          G    300.00   3500.00 1800.00      1
 1.12578097e+01 4.34354098e-02-2.02455774e-05 4.54245292e-09-4.01195170e-13    2
-2.30439963e+04-4.47863376e+01-9.43363126e+00 8.94163897e-02-5.85630607e-05    3
 1.87341134e-08-2.37225913e-12-1.55950776e+04 6.72000574e+01                   4
CYC6H8                  C   6H   8          G    300.00   3500.00 1490.00      1
 8.66772260e+00 3.45074855e-02-1.63846780e-05 3.69260975e-09-3.24421026e-13    2
 5.74022139e+03-2.73566208e+01-6.91358136e+00 7.63364895e-02-5.84944135e-05    3
 2.25336547e-08-3.48567018e-12 1.03834500e+04 5.40276160e+01                   4
CYC6H9                  C   6H   9          G    300.00   3500.00 1800.00      1
 1.41670463e+01 2.75651338e-02-1.13337615e-05 2.23021652e-09-1.74683445e-13    2
 7.93866332e+03-5.85441979e+01-6.48639356e+00 7.34616669e-02-4.95808724e-05    3
 1.63958131e-08-2.14212742e-12 1.53739017e+04 5.32365273e+01                   4
DCYC5                   C  10H  16          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748172e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
DECALIN                 C  10H  18          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748172e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
DIBZFUR                 C  12H   8O   1     G    300.00   3500.00 1410.00      1
 2.49525256e+01 3.24730728e-02-1.15459374e-05 1.79679054e-09-9.97833662e-14    2
-5.30753651e+03-1.13355893e+02-1.16970901e+01 1.36443614e-01-1.22152896e-04    3
 5.40932248e-08-9.37220078e-12 5.02765510e+03 7.60497478e+01                   4
DIFENET                 C  12H  10O   1     G    300.00   3500.00 1430.00      1
 1.71548107e+01 5.25374196e-02-2.45657222e-05 5.58244776e-09-4.99409896e-13    2
-3.29704394e+03-6.49985669e+01-8.57458099e+00 1.24507746e-01-1.00059071e-04    3
 4.07774824e-08-6.65238798e-12 4.06156207e+03 6.83336207e+01                   4
DIPE                    C   6H  14O   1     G    300.00   3500.00 1380.00      1
 1.11573928e+01 4.99175659e-02-2.25561386e-05 4.38444843e-09-3.06549364e-13    2
-4.59357929e+04-3.06117763e+01-2.50745274e+00 8.95258138e-02-6.56085820e-05    3
 2.51827303e-08-4.07435404e-12-4.21642955e+04 3.97144256e+01                   4
DME-OO                  C   2H   5O   3     G    300.00   3500.00  870.00      1
 3.58974575e+00 2.80960123e-02-1.49224205e-05 3.71355557e-09-3.53703711e-13    2
-1.93352293e+04 1.47278303e+01 5.41345468e+00 1.97111437e-02-4.65750394e-07    3
-7.36435253e-09 2.82960321e-12-1.96525546e+04 6.18346241e+00                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   3500.00 1800.00      1
 9.57989146e+00 2.53360331e-02-1.13706887e-05 2.45690684e-09-2.09295699e-13    2
-3.48199648e+04-1.16031904e+01 7.85487749e+00 2.91693975e-02-1.45651591e-05    3
 3.64004400e-09-3.73620304e-13-3.41989598e+04-2.26705495e+00                   4
DME-OQOOH               C   2H   4O   4     G    300.00   3500.00 1760.00      1
 1.54960865e+01 1.58758106e-03 2.24425901e-06-9.74237206e-10 1.03773065e-13    2
-4.69655432e+04-5.18401164e+01 3.62388957e+00 2.85698467e-02-2.07519902e-05    3
 7.73646324e-09-1.13354234e-12-4.27865299e+04 1.21478877e+01                   4
DME-QOOH                C   2H   5O   3     G    300.00   3500.00 1800.00      1
 9.52551493e+00 1.89562856e-02-9.27557330e-06 2.15192754e-09-1.93905680e-13    2
-1.72537528e+04-1.74698518e+01 5.12252607e+00 2.87407053e-02-1.74292564e-05    3
 5.17181016e-09-6.13333823e-13-1.56686768e+04 6.36004246e+00                   4
DMF                     C   6H   8O   1     G    300.00   3500.00 1590.00      1
 1.38889506e+01 2.49736923e-02-8.98421021e-06 1.42738238e-09-7.97717945e-14    2
-2.20872034e+04-4.94041109e+01-2.31533181e+00 6.57391826e-02-4.74422199e-05    3
 1.75523340e-08-2.61514155e-12-1.69342416e+04 3.62866615e+01                   4
DMF-3YL                 C   6H   7O   1     G    300.00   3500.00 1620.00      1
 1.41703395e+01 2.18230092e-02-7.69511407e-06 1.17891300e-09-6.12376638e-14    2
 1.19557792e+04-4.86583489e+01-1.12307984e+00 5.95845385e-02-4.26594930e-05    3
 1.55675463e-08-2.28170577e-12 1.69108471e+04 3.25015043e+01                   4
ERC4H8CHO               C   5H   9O   1     G    300.00   3500.00  750.00      1
-3.04813054e-01 5.67977502e-02-3.24057642e-05 8.50471985e-09-8.41763290e-13    2
-5.21420511e+03 3.41933259e+01 6.22525332e+00 2.19707295e-02 3.72482771e-05    3
-5.34099835e-08 1.97964712e-11-6.19371507e+03 4.56811339e+00                   4
ETBE                    C   6H  14O   1     G    300.00   3500.00 1280.00      1
 1.16559136e+01 4.67933987e-02-1.93342014e-05 3.59185140e-09-2.45564975e-13    2
-4.60322114e+04-3.38084939e+01-3.48005604e+00 9.40933039e-02-7.47637778e-05    3
 3.24614225e-08-5.88415307e-12-4.21574031e+04 4.29502770e+01                   4
ETC3H4O2                C   3H   4O   2     G    300.00   3500.00 1240.00      1
 1.02920429e+01 1.38871300e-02-6.12561993e-06 1.30548845e-09-1.09965765e-13    2
-3.57026988e+04-2.69350036e+01 1.17378045e-01 4.67086294e-02-4.58290467e-05    3
 2.26514168e-08-4.41358036e-12-3.31793820e+04 2.43405589e+01                   4
ETEROMD                 C  11H  20O   3     G    300.00   3500.00 1760.00      1
 4.14249213e+01 4.51122053e-02-1.56530088e-05 2.49214075e-09-1.50324737e-13    2
-8.95581279e+04-1.84296546e+02-1.24327962e-01 1.39542317e-01-9.61332178e-05    3
 3.29770684e-08-4.48057014e-12-7.49327921e+04 3.96429285e+01                   4
ETEROMPA                C  17H  32O   3     G    300.00   3500.00 1310.00      1
 4.32126695e+01 9.17256499e-02-3.02788098e-05 4.53882493e-09-2.50045022e-13    2
-1.06117741e+05-1.75617618e+02-8.73011664e+00 2.50329577e-01-2.11886360e-04    3
 9.69599701e-08-1.78876681e-11-9.25087311e+04 8.90022613e+01                   4
ETMB583                 C   5H   8O   3     G    300.00   3500.00 1270.00      1
 1.75630365e+01 2.35383857e-02-7.56913166e-06 1.05837457e-09-4.95698273e-14    2
-6.27369638e+04-6.15054259e+01-4.60165685e+00 9.33484435e-02-9.00219559e-05    3
 4.43406970e-08-8.56971204e-12-5.71071317e+04 5.07241435e+01                   4
FLUORENE                C  13H  10          G    300.00   3500.00 1440.00      1
 2.91248872e+01 2.85362024e-02-5.66199729e-06-5.67026725e-10 1.91134972e-13    2
 9.75119358e+03-1.37159218e+02-1.43465120e+01 1.49290089e-01-1.31447296e-04    3
 5.76669078e-08-9.91892310e-12 2.22709565e+04 8.84167006e+01                   4
GLIET                   C   2H   6O   2     G    300.00   3500.00 1470.00      1
 6.66621468e+00 1.87459315e-02-7.66039208e-06 1.53874843e-09-1.24203245e-13    2
-4.95959120e+04-6.01671900e+00 9.46220545e-01 3.43105414e-02-2.35426471e-05    3
 8.74158516e-09-1.34917548e-12-4.79142337e+04 2.37826449e+01                   4
GLYCEROL                C   3H   8O   3     G    300.00   3500.00 1290.00      1
 1.14796489e+01 2.36292461e-02-8.98384419e-06 1.70355137e-09-1.31527258e-13    2
-7.41781076e+04-2.56707288e+01 1.97850806e-01 5.86115658e-02-4.96609601e-05    3
 2.27253167e-08-4.20551279e-12-7.12674037e+04 3.16302477e+01                   4
H                       H   1               G    300.00   3500.00 1490.00      1
 2.50000000e+00 7.40336223e-15-5.56967416e-18 1.73924876e-21-1.92673709e-25    2
 2.54716200e+04-4.60117600e-01 2.50000000e+00-4.07455160e-15 5.98527266e-18    3
-3.43074982e-21 6.74775716e-25 2.54716200e+04-4.60117600e-01                   4
H2                      H   2               G    300.00   3500.00  750.00      1
 3.73110902e+00-8.86706214e-04 1.12286897e-06-3.74349782e-10 4.17963674e-14    2
-1.08851547e+03-5.35285855e+00 3.08866003e+00 2.53968841e-03-5.72992027e-06    3
 5.71701843e-09-1.98865970e-12-9.92148124e+02-2.43823459e+00                   4
H2CN                    C   1H   2N   1     G    300.00   3500.00 1800.00      1
 5.22111320e+00 3.42647499e-03-8.36137799e-07 4.74833030e-11 4.28153350e-15    2
 2.75312364e+04-4.80262216e+00 1.81354567e+00 1.09988473e-02-7.14644805e-06    3
 2.38463525e-09-3.20322903e-13 2.87579607e+04 1.36398442e+01                   4
H2NO                    H   2O   1N   1     G    300.00   3500.00 1200.00      1
 1.43405821e+00 9.01333883e-03-3.38828321e-06 4.28655869e-10-2.36936075e-15    2
 7.27341661e+03 1.79341864e+01 2.78935895e+00 4.49566971e-03 2.25880318e-06    3
-2.70861435e-09 6.51228601e-13 6.94814443e+03 1.11485432e+01                   4
H2O                     H   2O   1          G    300.00   3500.00 1590.00      1
 2.30940463e+00 3.65433887e-03-1.22983871e-06 2.11931683e-10-1.50333493e-14    2
-2.97294901e+04 8.92765177e+00 4.03530937e+00-6.87559833e-04 2.86629214e-06    3
-1.50552360e-09 2.55006790e-13-3.02783278e+04-1.99201641e-01                   4
H2O2                    H   2O   2          G    300.00   3500.00 1180.00      1
 4.56163072e+00 4.35560969e-03-1.48694629e-06 2.38275424e-10-1.46610352e-14    2
-1.80016693e+04 5.66597119e-01 2.91896355e+00 9.92397296e-03-8.56537418e-06    3
 4.23738723e-09-8.61930485e-13-1.76139998e+04 8.76340177e+00                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1800.00      1
 7.44900312e+00 1.01177830e-03 3.02918165e-07-2.13909391e-10 2.81815208e-14    2
 1.86458955e+04-1.30987733e+01 4.44514163e+00 7.68702606e-03-5.25978830e-06    3
 1.84635226e-09-2.57965931e-13 1.97272856e+04 3.15875175e+00                   4
HCN                     C   1H   1N   1     G    300.00   3500.00  850.00      1
 3.48152100e+00 3.81748410e-03-1.53642929e-06 3.02291150e-10-2.35861473e-14    2
 1.50427831e+04 3.30702298e+00 2.53139665e+00 8.28865751e-03-9.42673531e-06    3
 6.49076646e-09-1.84372594e-12 1.52043042e+04 7.73641055e+00                   4
HCNO                    C   1H   1O   1N   1G    300.00   3500.00 1350.00      1
 7.12423974e+00 1.61853378e-03 2.31339437e-07-2.53211924e-10 3.63453797e-14    2
 1.67567928e+04-1.48886865e+01 2.20954024e+00 1.61806064e-02-1.59487412e-05    3
 7.73695136e-09-1.44331449e-12 1.80837616e+04 1.02968215e+01                   4
HCO                     C   1H   1O   1     G    300.00   3500.00  920.00      1
 2.44772078e+00 5.65570555e-03-3.01329556e-06 7.57702524e-10-7.26129631e-14    2
 4.31149160e+03 1.15871953e+01 3.74218864e+00 2.75844059e-05 6.16298892e-06    3
-5.89177898e-09 1.73431136e-12 4.07330951e+03 5.45007090e+00                   4
HCO3                    C   1H   1O   3     G    300.00   3500.00 1800.00      1
 5.04067718e+00 8.66656109e-03-4.28958277e-06 1.00563376e-09-9.13599886e-14    2
-1.77902136e+04 5.78191516e+00 3.79300672e+00 1.14391621e-02-6.60008362e-06    3
 1.86137482e-09-2.10212913e-13-1.73410522e+04 1.25345680e+01                   4
HCO3H                   C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230668e+01 4.43563253e-03-1.56188514e-06 2.43424395e-10-1.38391379e-14    2
-3.81313332e+04-2.33590722e+01 2.47434199e+00 2.16898607e-02-1.63512235e-05    3
 5.87745807e-09-8.18701091e-13-3.54892796e+04 1.72835470e+01                   4
HCOOH                   C   1H   2O   2     G    300.00   3500.00 1800.00      1
 5.80573302e+00 6.82017393e-03-2.95480608e-06 6.14340060e-10-5.06753135e-14    2
-4.80534416e+04-6.42993389e+00 1.36256505e+00 1.66938805e-02-1.11828949e-05    3
 3.66178037e-09-4.73930912e-13-4.64539011e+04 1.76174180e+01                   4
HE                      HE  1               G    300.00   3500.00 1490.00      1
 2.50000000e+00 7.40336223e-15-5.56967416e-18 1.73924876e-21-1.92673709e-25    2
-7.45375000e+02 9.28723974e-01 2.50000000e+00-4.07455160e-15 5.98527266e-18    3
-3.43074982e-21 6.74775716e-25-7.45375000e+02 9.28723974e-01                   4
HNCO                    C   1H   1O   1N   1G    300.00   3500.00 1660.00      1
 7.29502452e+00 4.88032844e-04 8.74568316e-07-4.09105701e-10 5.01959355e-14    2
-1.52722297e+04-1.41696888e+01 2.99127956e+00 1.08585026e-02-8.49633812e-06    3
 3.35431054e-09-5.16583618e-13-1.38433864e+04 8.77460657e+00                   4
HNNO                    H   1O   1N   2     G    300.00   3500.00 1360.00      1
 4.88500308e+00 5.60936901e-03-2.60717829e-06 5.93839036e-10-5.41495114e-14    2
 2.58926738e+04 6.01980007e-01 2.29344827e+00 1.32315890e-02-1.10140386e-05    3
 4.71484900e-09-8.11688108e-13 2.65975767e+04 1.39015974e+01                   4
HNO                     H   1O   1N   1     G    300.00   3500.00  900.00      1
 2.72673666e+00 5.06770488e-03-2.61122761e-06 6.38493559e-10-6.01581004e-14    2
 1.09769405e+04 9.63912842e+00 3.40204752e+00 2.06632330e-03 2.39107502e-06    3
-3.06691580e-09 9.69122277e-13 1.08553846e+04 6.45229501e+00                   4
HNO2                    H   1O   2N   1     G    300.00   3500.00 1800.00      1
 3.30359406e+00 7.74006618e-03-3.91474332e-06 9.47112178e-10-8.88494507e-14    2
-8.65702544e+03 7.10072496e+00 1.68890715e+00 1.13282593e-02-6.90490427e-06    3
 2.05457920e-09-2.42664314e-13-8.07573815e+03 1.58397474e+01                   4
HO2                     H   1O   2          G    300.00   3500.00 1540.00      1
 4.16318067e+00 1.99798265e-03-4.89192086e-07 7.71153172e-11-7.30772104e-15    2
 4.41348948e+01 2.95517985e+00 2.85241381e+00 5.40257188e-03-3.80535043e-06    3
 1.51268170e-09-2.40354212e-13 4.47851086e+02 9.84483831e+00                   4
HOCN                    C   1H   1O   1N   1G    300.00   3500.00 1760.00      1
 6.92286755e+00 1.77083687e-04 1.06417841e-06-4.55819441e-10 5.43563991e-14    2
-3.77375638e+03-1.08544042e+01 3.05788784e+00 8.96112848e-03-6.42222341e-06    3
 2.37993882e-09-3.48450172e-13-2.41328352e+03 9.97681509e+00                   4
HONO                    H   1O   2N   1     G    300.00   3500.00 1420.00      1
 5.88742112e+00 3.49329101e-03-1.17730803e-06 1.65569378e-10-6.87715202e-15    2
-1.14386309e+04-5.23866548e+00 2.37883184e+00 1.33766411e-02-1.16174666e-05    3
 5.06705227e-09-8.69814280e-13-1.04421916e+04 1.29185606e+01                   4
HONO2                   H   1O   3N   1     G    300.00   3500.00 1310.00      1
 5.20949091e+00 9.97123440e-03-5.50725421e-06 1.39250696e-09-1.33157469e-13    2
-1.74464288e+04-1.35430787e+00 8.85706040e-01 2.31736309e-02-2.06245022e-05    3
 9.08576291e-09-1.60133609e-12-1.63135971e+04 2.06729940e+01                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1420.00      1
 4.21122112e+01 1.11834123e-01-5.11978482e-05 1.12541459e-08-9.72533984e-13    2
-7.89343498e+04-1.80495570e+02-6.54289827e+00 2.48890769e-01-1.95975996e-04    3
 7.92251073e-08-1.29392525e-11-6.51162987e+04 7.12984570e+01                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1590.00      1
 5.03105902e+01 8.85535013e-02-3.63077668e-05 7.13747183e-09-5.56692148e-13    2
-1.01978074e+05-2.30341253e+02-5.93668664e+00 2.30056085e-01-1.69800770e-04    3
 6.31093809e-08-9.35730677e-12-8.40914402e+04 6.71031189e+01                   4
IC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1460.00      1
 4.22439745e+01 1.02589738e-01-4.54459633e-05 9.70909447e-09-8.19911243e-13    2
-6.26654622e+04-1.86283114e+02-7.79323360e+00 2.39677979e-01-1.86290047e-04    3
 7.40214614e-08-1.18323028e-11-4.80545975e+04 7.40533932e+01                   4
IC16H33                 C  16H  33          G    300.00   3500.00 1650.00      1
 5.11453588e+01 7.53296743e-02-2.79263242e-05 4.92908201e-09-3.44364401e-13    2
-5.61938874e+04-2.43048234e+02-8.95216175e+00 2.21020633e-01-1.60372651e-04    3
 5.84427492e-08-8.45249579e-12-3.63617056e+04 7.69829165e+01                   4
IC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1460.00      1
 3.94749769e+01 1.06211481e-01-4.74108472e-05 1.02029370e-08-8.67107397e-13    2
-6.81954459e+04-1.73182708e+02-7.55515778e+00 2.35061165e-01-1.79790660e-04    3
 7.06503399e-08-1.12176901e-11-5.44626465e+04 7.15084222e+01                   4
IC16H34                 C  16H  34          G    300.00   3500.00 1590.00      1
 4.72524600e+01 8.54680758e-02-3.36612723e-05 6.38202029e-09-4.82094887e-13    2
-7.78744143e+04-2.24182950e+02-9.93612250e+00 2.29338723e-01-1.69388298e-04    3
 6.32906266e-08-9.42998897e-12-5.96884450e+04 7.82391931e+01                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   3500.00 1370.00      1
 4.07769110e+01 1.15135971e-01-5.36319133e-05 1.19826916e-08-1.04989886e-12    2
-8.16821240e+04-1.74509322e+02-7.08781179e+00 2.54886986e-01-2.06643974e-04    3
 8.64411154e-08-1.46372025e-11-6.85671899e+04 7.14786263e+01                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   3500.00 1560.00      1
 5.03537527e+01 8.72534729e-02-3.55849544e-05 6.99643634e-09-5.47405935e-13    2
-6.86134004e+04-2.32227161e+02-7.33743336e+00 2.35179591e-01-1.77821606e-04    3
 6.77813303e-08-1.02885748e-11-5.06137504e+04 7.17539151e+01                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1220.00      1
 1.23035624e+01 2.79964883e-02-1.33482910e-05 3.03524083e-09-2.69271163e-13    2
-2.25784829e+04-2.78550798e+01 1.73143843e+00 6.26591900e-02-5.59663668e-05    3
 2.63238068e-08-5.04151829e-12-1.99988847e+04 2.52515831e+01                   4
IC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1270.00      1
 1.04498043e+01 2.29490980e-02-1.05757759e-05 2.34172678e-09-2.03669153e-13    2
-5.22299426e+03-2.40008692e+01-1.71110880e-01 5.64007993e-02-5.00856593e-05    3
 2.30818231e-08-4.28636527e-12-2.52528181e+03 2.97774852e+01                   4
IC3H5CHO                C   4H   6O   1     G    300.00   3500.00 1370.00      1
 8.96605760e+00 2.20962385e-02-1.00901145e-05 2.22139279e-09-1.91792264e-13    2
-1.79920102e+04-2.11939239e+01 6.92941977e-01 4.62513206e-02-3.65372847e-05    3
 1.50910620e-08-2.54027204e-12-1.57251765e+04 2.13235423e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1630.00      1
 8.48779790e+00 1.53259253e-02-4.76474417e-06 3.92065263e-10 2.47111520e-14    2
 5.50507422e+03-2.12719618e+01 2.73725246e-01 3.54831588e-02-2.33143455e-05    3
 7.97881429e-09-1.13890066e-12 8.18286190e+03 2.23694223e+01                   4
IC3H7CHO                C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.25375038e+01 2.06759832e-02-7.90606663e-06 1.44761601e-09-1.05776578e-13    2
-3.22363635e+04-4.10505202e+01-3.44732114e-01 4.93031741e-02-3.17620591e-05    3
 1.02831688e-08-1.33293668e-12-2.75987585e+04 2.86708279e+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1310.00      1
 6.28069615e+00 2.59370043e-02-1.05350747e-05 1.92921360e-09-1.30183993e-13    2
-3.63768639e+04-6.66341882e+00-3.00574060e-01 4.60324859e-02-3.35451681e-05    3
 1.36391848e-08-2.36491132e-12-3.46525711e+04 2.68645272e+01                   4
IC3H7OO                 C   3H   7O   2     G    300.00   3500.00 1260.00      1
 7.34738699e+00 2.68252330e-02-1.24179691e-05 2.76645854e-09-2.42147350e-13    2
-1.06484855e+04-8.92587196e+00 1.07341266e+00 4.67426118e-02-3.61291344e-05    3
 1.53120486e-08-2.73135173e-12-9.06744395e+03 2.27924165e+01                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1570.00      1
 1.51567879e+01 2.57227734e-02-1.11020451e-05 2.28943519e-09-1.86269530e-13    2
-4.30658407e+04-4.59845002e+01 9.69279340e-01 6.18692920e-02-4.56369355e-05    3
 1.69539322e-08-2.52138051e-12-3.86109630e+04 2.88616666e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955794e+00 3.23747266e-02-1.18655436e-05 1.37455178e-09 1.57073476e-14    2
-1.97025810e+04-6.34483422e+00-1.85965328e+00 5.58007940e-02-3.97537190e-05    3
 1.61302002e-08-2.91200067e-12-1.78430198e+04 3.09610166e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177121e+00 3.67769036e-02-1.77031336e-05 3.74786262e-09-2.92191280e-13    2
 1.31214242e+04 2.00120538e+01 3.86129991e+00 2.14653110e-02 1.51074220e-05    3
-2.75002856e-08 1.08678616e-11 1.27462902e+04 8.04059744e+00                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433967e+00 2.47722696e-02-1.05415828e-05 2.18152373e-09-1.80119594e-13    2
-6.21385768e+03-1.72949366e+01 7.17301598e-01 4.01434653e-02-2.33509125e-05    3
 6.92571993e-09-8.39035734e-13-3.72372397e+03 2.01415164e+01                   4
IC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.44537517e+01 2.20810695e-02-7.57959310e-06 1.19533670e-09-7.16167606e-14    2
-4.15822810e+04-5.13315495e+01-5.45479447e-01 5.54126942e-02-3.53559470e-05    3
 1.14828752e-08-1.50044155e-12-3.61825578e+04 2.98474183e+01                   4
IC4H9P                  C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880517e+00 2.55088283e-02-8.62221491e-06 8.09648923e-10 4.02033219e-14    2
 3.37759298e+03-1.61084037e+01-1.15582376e+00 5.10042938e-02-3.53657102e-05    3
 1.32774789e-08-2.13948724e-12 5.98437685e+03 3.11244820e+01                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   3500.00 1380.00      1
 8.54295826e+00 3.45220773e-02-1.59311943e-05 3.53852672e-09-3.08950056e-13    2
-1.29532173e+04-1.39825068e+01 7.00555201e-01 5.72536803e-02-4.06394585e-05    3
 1.54748862e-08-2.47133403e-12-1.07887140e+04 2.63784632e+01                   4
IC4H9T                  C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871688e+00 2.55264450e-02-8.65284050e-06 8.24419704e-10 3.80550653e-14    2
 8.35470581e+02-1.73299272e+01-1.29900233e+00 5.18342142e-02-3.68397360e-05    3
 1.42467509e-08-2.35878979e-12 3.41363196e+03 3.01901373e+01                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   3500.00 1260.00      1
 9.11667611e+00 3.41757258e-02-1.58797345e-05 3.54686464e-09-3.10976548e-13    2
-1.64591648e+04-1.96564028e+01 4.84069009e-01 6.15808277e-02-4.85048558e-05    3
 2.08088336e-08-3.73597039e-12-1.42837478e+04 2.39860330e+01                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1290.00      1
 1.30518446e+01 3.65484801e-02-1.74274782e-05 3.96741952e-09-3.52552034e-13    2
-2.47096139e+04-3.04334702e+01 1.64511788e+00 7.19181753e-02-5.85550308e-05    3
 2.52219686e-08-4.47165070e-12-2.17666784e+04 2.75020267e+01                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   3500.00 1350.00      1
 1.14809469e+01 3.08095616e-02-1.41939360e-05 3.14755455e-09-2.74422165e-13    2
-7.45268236e+03-2.80879239e+01-1.93281563e-01 6.53998681e-02-5.26276099e-05    3
 2.21271466e-08-3.78916143e-12-4.30064068e+03 3.17369695e+01                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1240.00      1
 1.39939782e+01 3.54845222e-02-1.68915059e-05 3.83671077e-09-3.40131614e-13    2
-2.83614519e+04-3.70531088e+01 1.55094393e+00 7.56233424e-02-6.54465303e-05    3
 2.99415626e-08-5.60320657e-12-2.52755794e+04 2.56539769e+01                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   3500.00 1270.00      1
 1.20890742e+01 3.03954175e-02-1.40883982e-05 3.13822121e-09-2.74437748e-13    2
-1.09705556e+04-3.28537329e+01-4.26302143e-01 6.98139255e-02-6.06456912e-05    3
 2.75777451e-08-5.08536764e-12-7.79165002e+03 3.05171096e+01                   4
IC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 2.13459841e+01 8.88367161e-03 1.59648418e-06-1.31808203e-09 1.74600856e-13    2
-1.26620076e+04-8.94699897e+01-1.59634535e+00 5.98666259e-02-4.08893110e-05    3
 1.44173977e-08-2.01088244e-12-4.40276906e+03 3.46986831e+01                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   3500.00 1710.00      1
 3.48314225e+01 3.98146097e-02-1.43978345e-05 2.42273589e-09-1.57988116e-13    2
-5.01227380e+04-1.45334518e+02 1.76391327e+00 1.17165508e-01-8.22495000e-05    3
 2.88756269e-08-4.02536985e-12-3.88136498e+04 3.19375985e+01                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   3500.00 1770.00      1
 3.33140926e+01 3.48304479e-02-1.19632189e-05 1.85711682e-09-1.07309433e-13    2
-6.88276671e+04-1.40834098e+02 5.55148980e-01 1.08861959e-01-7.47017874e-05    3
 2.54874628e-08-3.44492892e-12-5.72310011e+04 3.59135548e+01                   4
IC8-QOOH                C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202581e+01 4.65574275e-02-1.91478836e-05 3.78861311e-09-2.97862012e-13    2
-2.91331926e+04-1.00455337e+02-9.92411236e-01 1.15564272e-01-8.55006187e-05    3
 3.21444828e-08-4.84207190e-12-2.07364398e+04 4.13504180e+01                   4
IC8H16                  C   8H  16          G    300.00   3500.00 1400.00      1
 1.88616063e+01 4.14292819e-02-1.28170544e-05 1.66806736e-09-6.58961711e-14    2
-2.24684067e+04-7.38514296e+01-5.35586581e+00 1.10622059e-01-8.69521729e-05    3
 3.69705048e-08-6.36990285e-12-1.56875145e+04 5.11323811e+01                   4
IC8H16O                 C   8H  16O   1     G    300.00   3500.00 1730.00      1
 2.92525449e+01 3.42835226e-02-1.16024061e-05 1.77291874e-09-1.00401812e-13    2
-4.92824114e+04-1.33818841e+02-8.05235857e+00 1.20537635e-01-8.63892084e-05    3
 3.05924957e-08-4.26508057e-12-3.63749148e+04 6.66033697e+01                   4
IC8H17                  C   8H  17          G    300.00   3500.00 1530.00      1
 2.65104230e+01 3.01796816e-02-5.82184991e-06 1.42085860e-11 7.60110759e-14    2
-1.80373025e+04-1.14981197e+02-3.32961207e+00 1.08192845e-01-8.23053435e-05    3
 3.33403496e-08-5.36943680e-12-8.90625182e+03 4.16697269e+01                   4
IC8H17-OO               C   8H  17O   2     G    300.00   3500.00 1600.00      1
 2.43863221e+01 4.79091863e-02-1.96116165e-05 3.85759153e-09-3.01446048e-13    2
-3.51809040e+04-9.31491997e+01-7.10506923e-01 1.10651259e-01-7.84323095e-05    3
 2.83662136e-08-4.13091825e-12-2.71499187e+04 3.97240936e+01                   4
IC8H18                  C   8H  18          G    300.00   3500.00 1390.00      1
 2.06155885e+01 4.43694094e-02-1.35968858e-05 1.75327622e-09-6.83090880e-14    2
-3.76580614e+04-8.42148793e+01-5.96912081e+00 1.20872170e-01-9.61538217e-05    3
 4.13489289e-08-7.18982936e-12-3.02675122e+04 5.27954202e+01                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202581e+01 4.65574275e-02-1.91478836e-05 3.78861311e-09-2.97862012e-13    2
-2.91331926e+04-1.00455337e+02-9.92411236e-01 1.15564272e-01-8.55006187e-05    3
 3.21444828e-08-4.84207190e-12-2.07364398e+04 4.13504180e+01                   4
INDENE                  C   9H   8          G    300.00   3500.00 1450.00      1
 1.65348693e+01 2.81361431e-02-7.82674558e-06 2.33936401e-10 1.15234436e-13    2
 1.13278665e+04-6.66478053e+01-7.32592199e+00 9.39590155e-02-7.59193723e-05    3
 3.15408912e-08-5.28251639e-12 1.82474960e+04 5.73325203e+01                   4
INDENYL                 C   9H   7          G    300.00   3500.00 1600.00      1
 1.63412613e+01 3.01210631e-02-1.29067938e-05 2.63187626e-09-2.11554314e-13    2
 2.91054096e+04-6.81510017e+01-5.81714820e+00 8.55170869e-02-6.48405661e-05    3
 2.42709481e-08-3.59265929e-12 3.61961007e+04 4.91650485e+01                   4
KEA3B3                  C   3H   4O   4     G    300.00   3500.00 1500.00      1
 1.56495498e+01 1.47904715e-02-6.84032429e-06 1.49167145e-09-1.26830372e-13    2
-4.74213138e+04-4.92482738e+01 1.41905665e+00 5.27384532e-02-4.47883060e-05    3
 1.83574411e-08-2.93779198e-12-4.31521659e+04 2.51755980e+01                   4
KEA3G2                  C   3H   4O   4     G    300.00   3500.00 1540.00      1
 1.52972938e+01 1.47507483e-02-6.65907582e-06 1.42291765e-09-1.19027510e-13    2
-5.03228961e+04-4.71892678e+01 2.76516864e+00 4.73017226e-02-3.83645703e-05    3
 1.51482399e-08-2.34716424e-12-4.64630015e+04 1.86821429e+01                   4
KEHYBU1                 C   4H   8O   4     G    300.00   3500.00 1200.00      1
 1.50812003e+01 2.99746636e-02-1.37944087e-05 3.03171375e-09-2.60935208e-13    2
-6.34178095e+04-4.27051069e+01-4.53521777e+00 9.53627237e-02-9.55294839e-05    3
 4.84400888e-08-9.72101335e-12-5.87098692e+04 5.55092666e+01                   4
KEHYMB                  C   5H   8O   5     G    300.00   3500.00 1200.00      1
 1.28585854e+01 3.05267697e-02-1.05263784e-05 1.70287735e-09-1.06411281e-13    2
-6.04915273e+04-3.42459469e+01-2.28352158e+00 8.10004596e-02-7.36184908e-05    3
 3.67540509e-08-7.40873910e-12-5.68574216e+04 4.15666988e+01                   4
KHDECA                  C  10H  16O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415883e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.98532958e+01-8.02402159e+00 8.95009509e-02-6.86853396e-05    3
 2.77298318e-08-4.50893790e-12-3.06512867e+04 5.22593733e+01                   4
KHMLIN1                 C  19H  30O   5     G    300.00   3500.00 1690.00      1
 6.18941987e+01 8.22994739e-02-3.10180668e-05 5.38913026e-09-3.62606874e-13    2
-9.79974660e+04-2.72277500e+02-3.09268744e+00 2.36114589e-01-1.67540358e-04    3
 5.92440776e-08-8.32931507e-12-7.60318984e+04 7.53471329e+01                   4
LC6H5                   C   6H   5          G    300.00   3500.00 1140.00      1
 1.23076076e+01 1.68261952e-02-6.51181371e-06 1.21158891e-09-8.99428218e-14    2
 5.89425072e+04-3.55373248e+01 1.67614175e-01 5.94226632e-02-6.25597980e-05    3
 3.39881879e-08-7.27779348e-12 6.17104257e+04 2.46218079e+01                   4
LC6H6                   C   6H   6          G    300.00   3500.00 1250.00      1
 1.28863876e+01 1.90072461e-02-7.30992558e-06 1.31482495e-09-9.21385789e-14    2
 3.55364843e+04-4.09021933e+01-1.05889383e+00 6.36321466e-02-6.08598062e-05    3
 2.98747613e-08-5.80412585e-12 3.90228046e+04 2.94875281e+01                   4
MACRIL                  C   4H   6O   2     G    300.00   3500.00 1110.00      1
 9.14034166e+00 2.10870489e-02-7.42259222e-06 1.25044332e-09-8.33064060e-14    2
-4.12827789e+04-1.50267978e+01-1.13135763e+00 5.81021815e-02-5.74430417e-05    3
 3.12927553e-08-6.84959289e-12-3.90024617e+04 3.56001684e+01                   4
MB                      C   5H  10O   2     G    300.00   3500.00 1800.00      1
 1.24284224e+01 3.57133446e-02-1.61592883e-05 3.52094113e-09-3.02693515e-13    2
-6.07702348e+04-3.65220690e+01 2.77831320e+00 5.71580318e-02-3.40298609e-05    3
 1.01396717e-08-1.22196165e-12-5.72961955e+04 1.57063351e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1540.00      1
 1.14154101e+01 2.70830264e-02-1.13419491e-05 2.30157826e-09-1.86056675e-13    2
 6.23040748e+03-4.10347479e+01-6.52219774e+00 7.36742157e-02-5.67229776e-05    3
 2.19470452e-08-3.37525585e-12 1.17551907e+04 5.32489849e+01                   4
MCROT                   C   5H   8O   2     G    300.00   3500.00 1270.00      1
 1.13738847e+01 2.61318034e-02-8.74855171e-06 1.35831508e-09-8.00175020e-14    2
-4.63062146e+04-2.54801461e+01 2.72064727e-01 6.10981657e-02-5.00474047e-05    3
 2.30375030e-08-4.34757418e-12-4.34863523e+04 3.07332406e+01                   4
MCYC6                   C   7H  14          G    300.00   3500.00 1800.00      1
 1.67194568e+01 4.36180644e-02-1.87773363e-05 3.92059023e-09-3.26702984e-13    2
-2.91866300e+04-7.40611877e+01-1.01006358e+01 1.03218270e-01-6.84441744e-05    3
 2.23157154e-08-2.88158149e-12-1.95313967e+04 7.10947481e+01                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587613e+01 3.12961497e-02-1.06604211e-05 1.62769455e-09-9.15073605e-14    2
-4.08526671e+04-1.40718316e+02-4.29317081e+00 1.12091476e-01-7.91310369e-05    3
 2.74170037e-08-3.73406515e-12-2.81964832e+04 5.21777121e+01                   4
MCYC6-OQOOH             C   7H  12O   3     G    300.00   3500.00 1800.00      1
 2.89245833e+01 2.89702632e-02-1.00807411e-05 1.60861341e-09-9.81376976e-14    2
-5.92858085e+04-1.29605491e+02-5.14358533e+00 1.04677305e-01-7.31699422e-05    3
 2.49749842e-08-3.34346697e-12-4.70212678e+04 5.47785441e+01                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659891e+01 2.65374271e-02-8.30522001e-06 1.12153176e-09-5.23348938e-14    2
-2.28599204e+04-1.33867706e+02-7.82169678e+00 1.09176729e-01-7.71713049e-05    3
 2.66274891e-08-3.59482897e-12-9.47235352e+03 6.73998075e+01                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587613e+01 3.12961497e-02-1.06604211e-05 1.62769455e-09-9.15073605e-14    2
-4.08526671e+04-1.40718316e+02-4.29317081e+00 1.12091476e-01-7.91310369e-05    3
 2.74170037e-08-3.73406515e-12-2.81964832e+04 5.21777121e+01                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659891e+01 2.65374271e-02-8.30522001e-06 1.12153176e-09-5.23348938e-14    2
-2.28599204e+04-1.33867706e+02-7.82169678e+00 1.09176729e-01-7.71713049e-05    3
 2.66274891e-08-3.59482897e-12-9.47235352e+03 6.73998075e+01                   4
MD                      C  11H  22O   2     G    300.00   3500.00 1800.00      1
 3.32942906e+01 6.02278032e-02-2.43433721e-05 4.77523421e-09-3.75629873e-13    2
-8.61538195e+04-1.40508531e+02 1.40263274e+00 1.31098154e-01-8.34019977e-05    3
 2.66487992e-08-3.41362502e-12-7.46728226e+04 3.20957740e+01                   4
MDKETO                  C  11H  20O   5     G    300.00   3500.00 1420.00      1
 2.98411867e+01 7.16595718e-02-3.12595573e-05 6.71204593e-09-5.73522120e-13    2
-1.08207342e+05-1.07784039e+02 3.72296254e+00 1.45232034e-01-1.08976947e-04    3
 4.31990835e-08-6.99729634e-12-1.00789766e+05 2.73798301e+01                   4
MEFU2                   C   5H   6O   1     G    300.00   3500.00 1260.00      1
 5.16398169e+00 3.29529080e-02-1.68209195e-05 4.03716052e-09-3.55511369e-13    2
-1.31841670e+04-2.67616710e+00-3.74149804e+00 6.12242723e-02-5.04773055e-05    3
 2.18447722e-08-3.88876765e-12-1.09399861e+04 4.23457855e+01                   4
MEK                     C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.00996674e+01 2.22850926e-02-8.24112797e-06 1.42760366e-09-9.77654881e-14    2
-3.40270944e+04-2.55002808e+01 1.67138626e+00 4.10146063e-02-2.38490560e-05    3
 7.20831776e-09-9.00642446e-13-3.09929132e+04 2.01153350e+01                   4
MEOLE                   C  19H  36O   2     G    300.00   3500.00 1800.00      1
 5.99431010e+01 8.58698597e-02-2.97675970e-05 4.64267973e-09-2.70021412e-13    2
-1.05323856e+05-2.71321378e+02-2.40342610e-02 2.19130160e-01-1.40817847e-04    3
 4.57724021e-08-5.98248285e-12-8.37356873e+04 5.32332675e+01                   4
MLIN1                   C  19H  32O   2     G    300.00   3500.00 1790.00      1
 6.02396272e+01 7.58944997e-02-2.57645248e-05 3.83449043e-09-2.03418185e-13    2
-7.74468689e+04-2.75096818e+02-2.53501097e+00 2.16173021e-01-1.43316358e-04    3
 4.76154339e-08-6.31807509e-12-5.49735485e+04 6.43028989e+01                   4
MLINO                   C  19H  34O   2     G    300.00   3500.00 1800.00      1
 6.05955674e+01 8.00185064e-02-2.72219227e-05 4.09057977e-09-2.22036540e-13    2
-9.16175365e+04-2.76065905e+02-1.22142744e+00 2.17389606e-01-1.41697839e-04    3
 4.64890673e-08-6.11071537e-12-6.93634183e+04 5.85005668e+01                   4
MPA                     C  17H  34O   2     G    300.00   3500.00 1570.00      1
 4.76347765e+01 8.91363271e-02-3.14080949e-05 4.73916072e-09-2.33379401e-13    2
-1.08404908e+05-2.13800451e+02-6.71212905e+00 2.27599781e-01-1.63698019e-04    3
 6.09132260e-08-9.17829426e-12-9.13399797e+04 7.29065166e+01                   4
MSTEA                   C  19H  38O   2     G    300.00   3500.00 1590.00      1
 5.57521885e+01 9.44092844e-02-3.21197984e-05 4.65296638e-09-2.12922185e-13    2
-1.17225837e+05-2.54579461e+02-7.52353560e+00 2.53593496e-01-1.82293583e-04    3
 6.76189138e-08-1.01132284e-11-9.71041567e+04 8.00324369e+01                   4
MSTEAKETO               C  19H  36O   5     G    300.00   3500.00 1630.00      1
 6.13348222e+01 9.80436966e-02-3.77033724e-05 6.80817282e-09-4.83388457e-13    2
-1.42870185e+05-2.70834349e+02-4.17722454e-01 2.49583683e-01-1.77157348e-04    3
 6.38445637e-08-9.23130116e-12-1.22738855e+05 5.72570421e+01                   4
MTBE                    C   5H  12O   1     G    300.00   3500.00 1320.00      1
 9.85250854e+00 4.01896195e-02-1.66704212e-05 3.10158953e-09-2.11537799e-13    2
-4.09274217e+04-2.61941109e+01-1.85856423e+00 7.56777188e-02-5.69978068e-05    3
 2.34689560e-08-4.06899357e-12-3.78356985e+04 3.35564110e+01                   4
MTBE-O                  C   5H  10O   2     G    300.00   3500.00 1520.00      1
 1.51388759e+01 2.99979380e-02-1.22799224e-05 2.46100800e-09-1.97690794e-13    2
-5.39879921e+04-5.57113238e+01-5.03717524e+00 8.30928094e-02-6.46761770e-05    3
 2.54418214e-08-3.97742985e-12-4.78544725e+04 5.00743811e+01                   4
MTBE-OO                 C   5H  11O   3     G    300.00   3500.00 1650.00      1
 1.64806404e+01 3.48147986e-02-1.47688716e-05 3.00165535e-09-2.41352124e-13    2
-3.59678540e+04-5.02874924e+01 2.84930352e+00 6.78604638e-02-4.48103854e-05    3
 1.51396407e-08-2.08044082e-12-3.14695128e+04 2.23020650e+01                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   3500.00 1360.00      1
 1.70053287e+01 4.31260455e-02-1.99573148e-05 4.44658587e-09-3.89314847e-13    2
-4.64302952e+04-4.61328184e+01 4.65469152e+00 7.94514489e-02-6.00220979e-05    3
 2.40861854e-08-3.99953536e-12-4.30709219e+04 1.72494984e+01                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   3500.00 1750.00      1
 2.60727575e+01 2.16561735e-02-7.50837024e-06 1.18094191e-09-6.95946679e-14    2
-6.60762157e+04-1.03020582e+02 2.39248713e+00 7.57825058e-02-5.39023694e-05    3
 1.88548464e-08-2.59443816e-12-5.77881211e+04 2.44748876e+01                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   3500.00 1320.00      1
 1.54436171e+01 3.66620452e-02-1.53964703e-05 3.18866664e-09-2.64826209e-13    2
-2.86187067e+04-4.25445321e+01 1.39866729e+00 7.92224991e-02-6.37606224e-05    3
 2.76150061e-08-4.89102686e-12-2.49108399e+04 2.91135557e+01                   4
N                       N   1               G    300.00   3500.00 1800.00      1
 2.43583682e+00 1.27743369e-04-8.58132365e-08 2.13268140e-11-1.23433516e-15    2
 5.61236145e+04 4.53259076e+00 2.50515554e+00-2.62982346e-05 4.25547663e-08    3
-2.62168907e-11 5.36895716e-15 5.60986597e+04 4.15742338e+00                   4
N1C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.19078661e+01 2.67959929e-02-1.07944841e-05 2.10106148e-09-1.63536607e-13    2
-3.95221179e+04-3.57389868e+01 7.73360084e-02 5.30860597e-02-3.27028730e-05    3
 1.02152796e-08-1.29051135e-12-3.52631271e+04 2.82903098e+01                   4
N2                      N   2               G    300.00   3500.00 1050.00      1
 2.71287897e+00 1.90359754e-03-8.54297556e-07 1.84170938e-10-1.54715988e-14    2
-8.40225273e+02 7.15926558e+00 3.85321336e+00-2.44053349e-03 5.35160392e-06    3
-3.75608397e-09 9.22684330e-13-1.07969550e+03 1.60217419e+00                   4
N2C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.39850075e+01 2.35768220e-02-8.73106106e-06 1.51546163e-09-1.02847459e-13    2
-4.24053999e+04-4.83702850e+01 1.11912948e-01 5.44059211e-02-3.44219770e-05    3
 1.10306157e-08-1.42439663e-12-3.74110858e+04 2.67137970e+01                   4
N2H2                    H   2N   2          G    300.00   3500.00  930.00      1
 1.94872574e+00 9.02206572e-03-4.48167913e-06 1.07159624e-09-9.96387287e-14    2
 2.46850174e+04 1.27074554e+01 2.44745784e+00 6.87698140e-03-1.02186571e-06    3
-1.40855675e-09 5.67069064e-13 2.45922533e+04 1.03375547e+01                   4
N2H3                    H   3N   2          G    300.00   3500.00 1610.00      1
 5.06961797e+00 6.18061831e-03-1.87909018e-06 2.33273638e-10-8.03110073e-15    2
 1.63477734e+04-4.00218491e+00 1.71415249e+00 1.45171785e-02-9.64607174e-06    3
 3.44941507e-09-5.07431944e-13 1.74282333e+04 1.37839838e+01                   4
N2H4                    H   4N   2          G    300.00   3500.00 1160.00      1
 4.91914378e+00 9.71187969e-03-3.62925367e-06 6.36530934e-10-4.28508947e-14    2
 9.36304606e+03-2.64395648e+00 3.60425651e-01 2.54315974e-02-2.39564748e-05    3
 1.23188419e-08-2.56059034e-12 1.04206687e+04 2.00258283e+01                   4
N2O                     O   1N   2          G    300.00   3500.00 1650.00      1
 5.52129143e+00 1.46645965e-03-3.04694075e-07-1.87106858e-11 8.50389041e-15    2
 7.81312268e+03-6.17451657e+00 2.68521969e+00 8.34178508e-03-6.55498992e-06    3
 2.50666137e-09-3.74128239e-13 8.74902635e+03 8.92812480e+00                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   3500.00 1800.00      1
 4.08087723e+01 4.96339543e-02-1.81420129e-05 3.12006732e-09-2.11175642e-13    2
-5.65432959e+04-1.73811020e+02 2.62701325e+00 1.34482308e-01-8.88489740e-05    3
 2.93078307e-08-3.84836500e-12-4.27978627e+04 3.28366249e+01                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   3500.00 1650.00      1
 2.99089271e+01 5.87016386e-02-2.37959516e-05 4.63914804e-09-3.59659107e-13    2
-7.07246459e+04-1.14602343e+02 2.87865509e+00 1.24229571e-01-8.33667990e-05    3
 2.87081773e-08-4.00648172e-12-6.18046561e+04 2.93391873e+01                   4
NC10-QOOH               C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.67714538e+01 4.56787199e-02-1.56929249e-05 2.49979255e-09-1.53467299e-13    2
-3.72897414e+04-1.54708984e+02 8.46533635e-01 1.25511876e-01-8.22205548e-05    3
 2.71396555e-08-3.57567048e-12-2.43567701e+04 3.97241784e+01                   4
NC10H19                 C  10H  19          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360661e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC10H20                 C  10H  20          G    300.00   3500.00 1800.00      1
 2.82971791e+01 4.89478938e-02-1.82737062e-05 3.23575201e-09-2.26811843e-13    2
-3.12534582e+04-1.16784058e+02-2.31417710e+00 1.16973130e-01-7.49614029e-05    3
 2.42311952e-08-3.14284562e-12-2.02333700e+04 4.88909878e+01                   4
NC10H21                 C  10H  21          G    300.00   3500.00 1800.00      1
 2.63212692e+01 5.52219738e-02-2.21266526e-05 4.33498891e-09-3.42316503e-13    2
-2.10175171e+04-1.03192977e+02-1.81057271e+00 1.17737178e-01-7.42226562e-05    3
 2.36298050e-08-3.02215208e-12-1.08900540e+04 4.90624204e+01                   4
NC10H21-OO              C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.23779830e+01 5.24885367e-02-1.93370131e-05 3.35369674e-09-2.28448799e-13    2
-4.06447276e+04-1.32098961e+02 1.67478189e+00 1.20717872e-01-7.61947929e-05    3
 2.44121337e-08-3.15323171e-12-2.95915752e+04 3.40731686e+01                   4
NC10H22                 C  10H  22          G    300.00   3500.00 1800.00      1
 2.92878918e+01 5.29920990e-02-1.98404553e-05 3.55616370e-09-2.54281184e-13    2
-4.56232379e+04-1.22752047e+02-2.17870143e+00 1.22917862e-01-7.81119243e-05    3
 2.51381893e-08-3.25178473e-12-3.42952643e+04 4.75517200e+01                   4
NC10MOOH                C  10H  20O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   3500.00 1800.00      1
 4.68889668e+01 5.84439691e-02-2.09491580e-05 3.49897609e-09-2.27324946e-13    2
-6.45487872e+04-2.03262107e+02 2.75932352e+00 1.56509843e-01-1.02670720e-04    3
 3.37662211e-08-4.43110898e-12-4.86621157e+04 3.55767286e+01                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   3500.00 1800.00      1
 2.89762540e+01 8.51935060e-02-4.32222039e-05 1.03184896e-08-9.52873634e-13    2
-7.66784457e+04-1.07151303e+02 4.95723376e+00 1.38569107e-01-8.77018710e-05    3
 2.67924404e-08-3.24092235e-12-6.80315984e+04 2.28446447e+01                   4
NC12-QOOH               C  12H  25O   2     G    300.00   3500.00 1800.00      1
 4.28763735e+01 5.51011626e-02-1.90602563e-05 3.05791504e-09-1.89217484e-13    2
-4.53973988e+04-1.84606456e+02 5.27389362e-01 1.49210016e-01-9.74843011e-05    3
 3.21038575e-08-4.22337617e-12-3.01517645e+04 4.45950809e+01                   4
NC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295229e-05 5.21804509e-09-4.10998518e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710595e-12-1.66984825e+04 5.11161660e+01                   4
NC12H25-OO              C  12H  25O   2     G    300.00   3500.00 1800.00      1
 3.82754174e+01 6.23046009e-02-2.29785783e-05 3.99220438e-09-2.72630412e-13    2
-4.86703034e+04-1.60846136e+02 1.39669302e+00 1.44257322e-01-9.12725124e-05    3
 2.92862540e-08-3.78569287e-12-3.53939626e+04 3.87492139e+01                   4
NC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414095e+01 6.11045883e-02-2.24641073e-05 3.93182440e-09-2.73349362e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1800.00      1
 5.83925916e+01 7.87490301e-02-2.86987240e-05 4.90944000e-09-3.29403315e-13    2
-8.05061539e+04-2.59209019e+02 2.14519035e+00 2.03743255e-01-1.32860578e-04    3
 4.34879045e-08-5.68752339e-12-6.02570894e+04 4.52136503e+01                   4
NC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1690.00      1
 4.88441297e+01 8.47833151e-02-3.17577492e-05 5.56702742e-09-3.82331487e-13    2
-9.50808904e+04-2.07202631e+02 1.75040694e+00 1.96247748e-01-1.30690678e-04    3
 4.45938236e-08-6.15552619e-12-7.91632121e+04 4.47087787e+01                   4
NC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.49634696e+01 7.74662171e-02-2.71265902e-05 4.36953904e-09-2.68719606e-13    2
-8.49949222e+04-2.46825964e+02 8.02842616e-02 1.99428851e-01-1.28762119e-04    3
 4.20123273e-08-5.49688464e-12-6.52369755e+04 5.02132837e+01                   4
NC16H33                 C  16H  33          G    300.00   3500.00 1800.00      1
 4.66278372e+01 8.00212238e-02-3.03236333e-05 5.55903616e-09-4.09822553e-13    2
-4.61545210e+04-2.04019481e+02-3.22413374e+00 1.90803381e-01-1.22642098e-04    3
 3.97510601e-08-5.15871477e-12-2.82078115e+04 6.57897858e+01                   4
NC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.00344484e+01 8.20070153e-02-3.03042993e-05 5.28016700e-09-3.62022840e-13    2
-6.47045872e+04-2.18137205e+02 8.65096715e-01 1.91272241e-01-1.21358654e-04    3
 3.90040022e-08-5.04588884e-12-4.70036206e+04 4.79775838e+01                   4
NC16H34                 C  16H  34          G    300.00   3500.00 1800.00      1
 4.98210237e+01 7.73881688e-02-2.77557896e-05 4.69678103e-09-3.12959243e-13    2
-7.08514664e+04-2.24842855e+02-3.64057977e+00 1.96191732e-01-1.26758759e-04    3
 4.13645475e-08-5.40570458e-12-5.16052891e+04 6.45024955e+01                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1260.00      1
 1.11683562e+01 2.95822139e-02-1.42526305e-05 3.27126849e-09-2.92476812e-13    2
-2.00281219e+04-2.06289848e+01 2.57588692e+00 5.68598942e-02-4.67260594e-05    3
 2.04529769e-08-3.70154594e-12-1.78628196e+04 2.28105329e+01                   4
NC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1800.00      1
 1.29748618e+01 1.76433870e-02-7.16935406e-06 1.42696153e-09-1.14477043e-13    2
-5.86411825e+03-3.67690498e+01 1.55643299e+00 4.30176732e-02-2.83145926e-05    3
 9.25853134e-09-1.20219507e-12-1.75348388e+03 2.50298688e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1650.00      1
 8.44692954e+00 1.52881013e-02-4.72394213e-06 3.72053769e-10 2.77825399e-14    2
 7.24499466e+03-1.97652064e+01 5.40130268e-01 3.44560996e-02-2.21493951e-05    3
 7.41264082e-09-1.03897307e-12 9.85423842e+03 2.23400592e+01                   4
NC3H7O                  C   3H   7O   1     G    300.00   3500.00 1800.00      1
 9.66226461e+00 1.80582994e-02-6.80752580e-06 1.22634214e-09-8.79552073e-14    2
-9.72942766e+03-2.55365895e+01-5.52121379e-01 4.07569349e-02-2.57230554e-05    3
 8.23209384e-09-1.06097628e-12-6.05224870e+03 2.97457983e+01                   4
NC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1800.00      1
 1.03578665e+01 1.87834500e-02-6.54155125e-06 1.06792692e-09-6.79101580e-14    2
-3.60054458e+04-2.89224528e+01 2.34636347e-01 4.12795171e-02-2.52882738e-05    3
 8.01115750e-09-1.03224774e-12-3.23610829e+04 2.58665808e+01                   4
NC3H7OO                 C   3H   7O   2     G    300.00   3500.00 1650.00      1
 9.25591855e+00 2.27563801e-02-9.54934453e-06 1.92559464e-09-1.53946670e-13    2
-9.34005086e+03-1.86388081e+01 1.92964396e+00 4.05170458e-02-2.56954042e-05    3
 8.44925513e-09-1.14238008e-12-6.92238025e+03 2.03750491e+01                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   3500.00 1230.00      1
 1.51474113e+01 3.37812811e-02-1.58996825e-05 3.57608795e-09-3.14486517e-13    2
-2.85698876e+04-4.24732203e+01 1.10123476e+00 7.94599040e-02-7.16053202e-05    3
 3.37688455e-08-6.45122586e-12-2.51145282e+04 2.81992197e+01                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1330.00      1
 1.18153445e+01 3.20093755e-02-1.53334981e-05 3.50316407e-09-3.12136547e-13    2
-4.27660549e+04-2.73083214e+01 2.51946600e+00 5.99669047e-02-4.68645461e-05    3
 1.93082006e-08-3.28300808e-12-4.02933512e+04 2.01899074e+01                   4
NC4-QOOH                C   4H   9O   2     G    300.00   3500.00 1760.00      1
 1.83774568e+01 1.83354725e-02-6.23923380e-06 9.66797421e-10-5.61281943e-14    2
-1.29135491e+04-6.55986639e+01 1.19976578e+00 5.73756794e-02-3.95121374e-05    3
 1.35701700e-08-1.84637998e-12-6.86700189e+03 2.69845517e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355362e+01 1.56272553e-02-3.14852000e-06-5.94424182e-11 5.32964635e-14    2
-2.28455262e+04-6.02417835e+01-1.20836758e+00 5.26137081e-02-3.39705640e-05    3
 1.13561294e-08-1.53219963e-12-1.68537208e+04 2.98384958e+01                   4
NC4H8                   C   4H   8          G    300.00   3500.00 1170.00      1
 2.98709814e+00 3.25282541e-02-1.46250479e-05 2.94136385e-09-2.14960813e-13    2
-2.50111901e+03 1.03971909e+01-1.05707773e+00 4.63544964e-02-3.23509995e-05    3
 1.30416212e-08-2.37313546e-12-1.55478186e+03 3.05429525e+01                   4
NC4H9-OO                C   4H   9O   2     G    300.00   3500.00 1320.00      1
 8.96630114e+00 3.41074657e-02-1.57641000e-05 3.50715782e-09-3.06662916e-13    2
-1.40847395e+04-1.58347447e+01 9.44281655e-01 5.84166156e-02-4.33881341e-05    3
 1.74586902e-08-2.94899859e-12-1.19669263e+04 2.50940293e+01                   4
NC4H9P                  C   4H   9          G    300.00   3500.00  950.00      1
 3.94763005e+00 3.16286394e-02-1.12984867e-05 1.11637452e-09 5.54031592e-14    2
 6.05554723e+03 7.76350069e+00-2.76188363e-01 4.94131380e-02-3.93792739e-05    3
 2.08221901e-08-5.13033778e-12 6.85807273e+03 2.79243294e+01                   4
NC4H9S                  C   4H   9          G    300.00   3500.00  850.00      1
 3.40122925e+00 3.20901864e-02-1.12255471e-05 9.71712129e-10 8.30726251e-14    2
 4.66283102e+03 1.05291640e+01 2.36336476e-01 4.69837994e-02-3.75083937e-05    3
 2.15857094e-08-5.97986776e-12 5.20086279e+03 2.52835872e+01                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   3500.00 1270.00      1
 1.54638476e+01 4.30531975e-02-2.04284728e-05 4.63174721e-09-4.10271992e-13    2
-3.17413365e+04-4.31406917e+01 1.43265566e+00 8.72459280e-02-7.26246113e-05    3
 3.20312950e-08-5.80388375e-12-2.81774138e+04 2.79053907e+01                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   3500.00 1410.00      1
 1.42172630e+01 3.77707683e-02-1.76257936e-05 3.93443034e-09-3.43954252e-13    2
-4.65061050e+04-3.85369191e+01 2.52749929e+00 7.09332187e-02-5.29049961e-05    3
 2.06149043e-08-3.30148510e-12-4.32095916e+04 2.18759162e+01                   4
NC5-QOOH                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.36538194e+01 3.77860020e-02-1.75151081e-05 3.90394425e-09-3.41708560e-13    2
-1.43879859e+04-3.94678819e+01-5.74283055e-01 8.15647789e-02-6.80290814e-05    3
 2.98085460e-08-5.32336273e-12-1.06886793e+04 3.29074336e+01                   4
NC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 1.11929736e+01 2.82582223e-02-1.13863841e-05 2.22526491e-09-1.74280993e-13    2
-1.02483443e+04-3.39253533e+01-6.89551964e-01 5.46638348e-02-3.33910611e-05    3
 1.03751453e-08-1.30620882e-12-5.97063504e+03 3.03853541e+01                   4
NC5H10-O                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.40073101e+01 3.04405284e-02-1.35854526e-05 2.90305354e-09-2.44985844e-13    2
-2.55455866e+04-5.25239383e+01-3.79263098e+00 6.99959530e-02-4.65483064e-05    3
 1.51115179e-08-1.94060590e-12-1.91376078e+04 4.38130562e+01                   4
NC5H11                  C   5H  11          G    300.00   3500.00 1800.00      1
 6.93193785e+00 3.75440987e-02-1.65478566e-05 3.53633643e-09-2.99976701e-13    2
-1.73087074e+03-8.88710670e+00-3.57520449e+00 6.08933039e-02-3.60055276e-05    3
 1.07428812e-08-1.30088570e-12 2.05170050e+03 4.79797395e+01                   4
NC5H11OOH               C   5H  12O   2     G    300.00   3500.00 1630.00      1
 1.66988185e+01 3.44172712e-02-1.43139761e-05 2.85300849e-09-2.25350876e-13    2
-3.73755763e+04-5.75775303e+01 6.24289371e-02 7.52427671e-02-5.18834508e-05    3
 1.82188468e-08-2.58207455e-12-3.19521133e+04 3.08116402e+01                   4
NC5H12                  C   5H  12          G    300.00   3500.00 1800.00      1
 2.12559082e+01 1.49866375e-02-1.56738312e-06-4.84518435e-10 9.00436509e-14    2
-2.80668702e+04-9.05497671e+01-1.97000865e+00 6.65997861e-02-4.45783403e-05    3
 1.54454657e-08-2.12245414e-12-1.97055401e+04 3.51537401e+01                   4
NC5H12OO                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.06544848e+01 4.16170555e-02-1.93382868e-05 4.32113942e-09-3.79088223e-13    2
-1.98652039e+04-2.50234586e+01 3.19664880e-01 7.34165014e-02-5.60299551e-05    3
 2.31373796e-08-3.99759595e-12-1.71781508e+04 2.75475609e+01                   4
NC5H9-3                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360661e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC6H12                  C   6H  12          G    300.00   3500.00 1780.00      1
 2.80951654e+01 5.24635942e-03 6.43208138e-06-3.19131389e-09 4.01093698e-13    2
-1.79767847e+04-1.24497292e+02-1.85358315e+00 7.25469181e-02-5.02818725e-05    3
 1.80498673e-08-2.58221827e-12-7.31503024e+03 3.72569567e+01                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   3500.00 1690.00      1
 2.24694069e+01 4.29307086e-02-1.68910162e-05 3.18431082e-09-2.38592446e-13    2
-4.58962940e+04-7.93472401e+01 2.87430503e+00 8.93096479e-02-5.80557552e-05    3
 1.94228666e-08-2.64074567e-12-3.92731495e+04 2.54699082e+01                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   3500.00 1670.00      1
 2.27584121e+01 4.25741258e-02-1.77950010e-05 3.55398722e-09-2.80791799e-13    2
-5.95329656e+04-8.19251639e+01 2.24997334e+00 9.16961348e-02-6.19165660e-05    3
 2.11673864e-08-2.91752820e-12-5.26831470e+04 2.75334100e+01                   4
NC7-QOOH                C   7H  15O   2     G    300.00   3500.00 1800.00      1
 3.67777501e+01 2.43465392e-02-1.65378817e-05 5.22869888e-09-5.85107382e-13    2
-2.84549794e+04-1.65059640e+02-2.87358792e+00 1.12460624e-01-8.99662853e-05    3
 3.24244039e-08-4.36228864e-12-1.41804977e+04 4.95416730e+01                   4
NC7H13                  C   7H  13          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360661e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC7H13OOH               C   7H  14O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC7H14                  C   7H  14          G    300.00   3500.00 1800.00      1
 1.82668105e+01 3.59607890e-02-1.37346402e-05 2.52229050e-09-1.85248240e-13    2
-1.87497345e+04-6.92309265e+01-1.22797309e+00 7.92825302e-02-4.98360912e-05    3
 1.58931983e-08-2.04231877e-12-1.17316124e+04 3.62789089e+01                   4
NC7H14O                 C   7H  14O   1     G    300.00   3500.00 1490.00      1
 1.37609323e+01 4.99379374e-02-2.21152348e-05 4.72010363e-09-3.98160014e-13    2
-3.97917916e+04-4.67908592e+01-7.39181743e+00 1.06723843e-01-7.92822536e-05    3
 3.02981881e-08-4.68978493e-12-3.34882722e+04 6.36941424e+01                   4
NC7H15                  C   7H  15          G    300.00   3500.00 1800.00      1
 1.58938298e+01 4.32851195e-02-1.83429598e-05 3.81524632e-09-3.18291961e-13    2
-8.33589206e+03-5.34387877e+01-1.03213606e+00 8.08983770e-02-4.96873411e-05    3
 1.54242764e-08-1.93065725e-12-2.24254435e+03 3.81680705e+01                   4
NC7H15-OO               C   7H  15O   2     G    300.00   3500.00 1780.00      1
 2.68006146e+01 3.35780866e-02-1.17982179e-05 1.89992229e-09-1.16218734e-13    2
-2.33388920e+04-1.06550436e+02 1.92333992e+00 8.94820746e-02-5.89083201e-05    3
 1.95441553e-08-2.59434135e-12-1.44825822e+04 2.78126029e+01                   4
NC7H15OOH               C   7H  16O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC7H16                  C   7H  16          G    300.00   3500.00 1800.00      1
 3.10696120e+01 1.73458864e-02-4.57663884e-07-1.06280964e-09 1.59098857e-13    2
-3.76541592e+04-1.40920497e+02-2.76912812e+00 9.25430866e-02-6.31219974e-05    3
 2.21462028e-08-3.06437509e-12-2.54722127e+04 4.22218230e+01                   4
NCO                     C   1O   1N   1     G    300.00   3500.00 1700.00      1
 5.80612871e+00 1.29457396e-03-2.96387145e-07-4.45669057e-12 6.00806513e-15    2
 1.70053704e+04-6.33800183e+00 2.87969597e+00 8.18029805e-03-6.37202605e-06    3
 2.37814680e-09-3.44374801e-13 1.80003575e+04 9.33319238e+00                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   3500.00 1800.00      1
 2.53088279e+01 2.46008468e-02-8.38584870e-06 1.28446216e-09-7.25492020e-14    2
-3.52662111e+04-9.88693150e+01 2.93992987e+00 7.43095092e-02-4.98097340e-05    3
 1.66266419e-08-2.20340750e-12-2.72134078e+04 2.21958278e+01                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   3500.00 1690.00      1
 2.24459936e+01 2.37621277e-02-8.83881473e-06 1.53830075e-09-1.04514815e-13    2
-5.03880249e+04-8.77405631e+01 1.27283562e+00 7.38761111e-02-5.33186817e-05    3
 1.90845993e-08-2.70012112e-12-4.32314975e+04 2.55178450e+01                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   3500.00 1630.00      1
 1.86197530e+01 2.85111424e-02-1.13969334e-05 2.18137254e-09-1.65768942e-13    2
-1.50391446e+04-6.74883738e+01 1.48070310e+00 7.05701605e-02-5.01015514e-05    3
 1.80114821e-08-2.59369986e-12-9.45181437e+03 2.35714319e+01                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   3500.00 1470.00      1
 1.29296103e+01 3.16150611e-02-1.35584975e-05 2.81753187e-09-2.32686285e-13    2
-2.37933924e+04-4.88968548e+01-6.91462638e+00 8.56129839e-02-6.86584188e-05    3
 2.78061583e-08-4.48245268e-12-1.79591868e+04 5.44853542e+01                   4
NEOC5H11                C   5H  11          G    300.00   3500.00 1670.00      1
 1.43276289e+01 2.66845577e-02-1.02158264e-05 1.86929104e-09-1.35803312e-13    2
-2.94216421e+03-5.15145769e+01-1.29689709e+00 6.41085720e-02-4.38302105e-05    3
 1.52882069e-08-2.14462305e-12 2.27642747e+03 3.18773552e+01                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   3500.00 1660.00      1
 1.69989732e+01 3.01601499e-02-1.19254896e-05 2.25822367e-09-1.69878947e-13    2
-2.10464569e+04-6.14617731e+01 1.07910948e+00 6.85212672e-02-4.65891499e-05    3
 1.61793724e-08-2.26643749e-12-1.57610621e+04 2.34108339e+01                   4
NEOC5H12                C   5H  12          G    300.00   3500.00 1700.00      1
 1.58220811e+01 2.73824077e-02-1.01392581e-05 1.77707009e-09-1.22756971e-13    2
-2.85197010e+04-6.62488521e+01-2.62463460e+00 7.07864446e-02-4.84369376e-05    3
 1.67957680e-08-2.33138901e-12-2.22478177e+04 3.25342362e+01                   4
NH                      H   1N   1          G    300.00   3500.00 1550.00      1
 2.53691464e+00 1.74532708e-03-6.66818142e-07 1.34160653e-10-1.04190033e-14    2
 4.21821879e+04 7.12732805e+00 3.75007687e+00-1.38541418e-03 2.36293147e-06    3
-1.16895746e-09 1.99761337e-13 4.18061076e+04 7.42847188e-01                   4
NH2                     H   2N   1          G    300.00   3500.00 1120.00      1
 2.67687765e+00 3.48484078e-03-1.28570820e-06 2.72091630e-10-2.36034281e-14    2
 2.20303372e+04 7.34730162e+00 4.18313061e+00-1.89463407e-03 5.91894562e-06    3
-4.01639279e-09 9.33647558e-13 2.16929365e+04-9.01998745e-02                   4
NH3                     H   3N   1          G    300.00   3500.00 1210.00      1
 2.21117984e+00 6.52182453e-03-2.30931532e-06 3.98907128e-10-2.80385645e-14    2
-6.39009604e+03 8.86905603e+00 3.21689186e+00 3.19715670e-03 1.81217371e-06    3
-1.87188573e-09 4.41133513e-13-6.63347835e+03 3.82536772e+00                   4
NNH                     H   1N   2          G    300.00   3500.00  720.00      1
 2.67540125e+00 5.35668680e-03-2.94990450e-06 7.78541240e-10-7.91413867e-14    2
 2.84746064e+04 1.03028707e+01 3.96823590e+00-1.82572793e-03 1.20134595e-05    3
-1.30764254e-08 4.73161093e-12 2.82884383e+04 4.49039228e+00                   4
NO                      O   1N   1          G    300.00   3500.00  970.00      1
 2.69775018e+00 2.39887133e-03-1.31644700e-06 3.38235813e-10-3.29394890e-14    2
 9.99854348e+03 9.40230813e+00 3.91290193e+00-2.61206371e-03 6.43242163e-06    3
-4.98744709e-09 1.33965920e-12 9.76280404e+03 3.57691592e+00                   4
NO2                     O   2N   1          G    300.00   3500.00 1800.00      1
 5.25673685e+00 1.64343307e-03-6.24197948e-07 1.07065150e-10-6.88584753e-15    2
 1.95363563e+03-2.35827568e+00 2.61409592e+00 7.51596848e-03-5.51797745e-06    3
 1.91957608e-09-2.58623476e-13 2.90498637e+03 1.19442483e+01                   4
NO3                     O   3N   1          G    300.00   3500.00 1330.00      1
 7.66391925e+00 2.28165967e-03-8.16241554e-07 1.11367864e-10-3.38429715e-15    2
 5.62975022e+03-1.51899442e+01 4.06541943e-01 2.41083583e-02-2.54328190e-05    3
 1.24505044e-08-2.32277087e-12 7.56021258e+03 2.18923574e+01                   4
NPBENZ                  C   9H  12          G    300.00   3500.00 1600.00      1
 1.88963371e+01 3.80090295e-02-1.52789389e-05 2.95630099e-09-2.27699217e-13    2
-8.96605283e+03-7.62711275e+01-5.58650157e+00 9.92161261e-02-7.26605920e-05    3
 2.68653231e-08-3.96348393e-12-1.13154446e+03 5.33514397e+01                   4
O                       O   1               G    300.00   3500.00  950.00      1
 2.57318360e+00-8.95609984e-05 4.05096303e-08-8.39812674e-12 9.43621991e-16    2
 2.92191409e+04 4.74952023e+00 2.95200330e+00-1.68459131e-03 2.55897854e-06    3
-1.77574473e-09 4.66034833e-13 2.91471652e+04 2.94136507e+00                   4
O2                      O   2               G    300.00   3500.00  760.00      1
 2.81750648e+00 2.49838007e-03-1.52493521e-06 4.50547608e-10-4.87702792e-14    2
-9.31713392e+02 7.94729337e+00 3.46035080e+00-8.85011121e-04 5.15281056e-06    3
-5.40712413e-09 1.87809542e-12-1.02942573e+03 5.02236126e+00                   4
ODECAL                  C  10H  18          G    300.00   3500.00 1800.00      1
 2.82109941e+01 4.74108396e-02-1.82963852e-05 3.42084161e-09-2.57817125e-13    2
-2.68355230e+04-1.31410203e+02-1.02710769e+01 1.32926553e-01-8.95594797e-05    3
 2.98145803e-08-3.92361417e-12-1.29819774e+04 7.68627930e+01                   4
OH                      H   1O   1          G    300.00   3500.00  880.00      1
 3.62538436e+00-5.02165281e-04 8.36958463e-07-2.95714531e-10 3.30350486e-14    2
 3.41380110e+03 1.55419440e+00 3.37995109e+00 6.13440526e-04-1.06464235e-06    3
 1.14489214e-09-3.76228211e-13 3.45699735e+03 2.70689352e+00                   4
PC3H4                   C   3H   4          G    300.00   3500.00  920.00      1
 3.04156590e+00 1.80732925e-02-9.19849468e-06 2.29161583e-09-2.25689445e-13    2
 2.06214251e+04 7.37493873e+00 1.35943188e+00 2.53869187e-02-2.11228852e-05    3
 1.09324785e-08-2.57374996e-12 2.09309378e+04 1.53500040e+01                   4
QBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1270.00      1
 9.44680463e+00 1.40890825e-02-6.70668585e-06 1.51288685e-09-1.32818576e-13    2
 1.91332917e+04-2.81812927e+01-5.88861871e+00 6.23896285e-02-6.37545748e-05    3
 3.14592852e-08-6.02777889e-12 2.30284892e+04 4.94686856e+01                   4
QDECOOH                 C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
QMBOOX                  C   5H   9O   4     G    300.00   3500.00 1350.00      1
 2.46557066e+01 1.60203243e-02-2.33018024e-06-2.09432791e-10 5.96256606e-14    2
-5.87318865e+04-9.28197844e+01-3.02577545e+00 9.80395304e-02-9.34626315e-05    3
 4.47942468e-08-8.27438909e-12-5.12578864e+04 4.90347050e+01                   4
QMDOOH                  C  11H  21O   4     G    300.00   3500.00 1800.00      1
 3.77681786e+01 6.05584838e-02-2.66377343e-05 5.63139231e-09-4.71383628e-13    2
-7.68263296e+04-1.55143375e+02 4.12866858e+00 1.35312950e-01-8.89331232e-05    3
 2.87037586e-08-3.67587894e-12-6.47161060e+04 2.69206708e+01                   4
QMEOLEOOH               C  19H  35O   4     G    300.00   3500.00 1800.00      1
 6.66288425e+01 8.44466273e-02-2.89700155e-05 4.40900507e-09-2.44932292e-13    2
-1.50877986e+05-3.00442019e+02-9.98790182e-01 2.34730256e-01-1.54206372e-04    3
 5.07928409e-08-6.68713172e-12-1.26532038e+05 6.55728373e+01                   4
QMLIN1OOX               C  19H  31O   4     G    300.00   3500.00 1610.00      1
 5.66825541e+01 9.03049166e-02-3.59434818e-05 6.72610917e-09-4.95506768e-13    2
-6.74923687e+04-2.44601780e+02-2.71828911e+00 2.37884651e-01-1.73440129e-04    3
 6.36605386e-08-9.33625668e-12-4.83652972e+04 7.02616632e+01                   4
QMLINOOX                C  19H  33O   4     G    300.00   3500.00 1760.00      1
 6.81309948e+01 7.45379902e-02-2.47878007e-05 3.55693559e-09-1.75307126e-13    2
-8.29474454e+04-3.08878538e+02 1.76458104e-02 2.29341056e-01-1.56722232e-04    3
 5.35320989e-08-7.27405191e-12-5.89715465e+04 5.82344142e+01                   4
QMPAOOH                 C  17H  33O   4     G    300.00   3500.00 1800.00      1
 3.77681786e+01 6.05584838e-02-2.66377343e-05 5.63139231e-09-4.71383628e-13    2
-7.68263296e+04-1.55143375e+02 4.12866858e+00 1.35312950e-01-8.89331232e-05    3
 2.87037586e-08-3.67587894e-12-6.47161060e+04 2.69206708e+01                   4
QMSTEAOOH               C  19H  37O   4     G    300.00   3500.00 1230.00      1
-1.30612117e+02 6.00365422e-01-4.85197519e-04 1.58690698e-07-1.80918283e-11    2
 1.24045727e+04 7.12083761e+02 2.15554530e+01 1.05511535e-01 1.18282831e-04    3
-1.68398923e-07 4.83898018e-11-2.50286496e+04-5.35376470e+01                   4
RALD3B                  C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013768e+00 4.60180077e-02-2.61696720e-05 6.65382129e-09-6.35305356e-13    2
-2.14966002e+03 5.90959839e+01 7.04072885e+00-2.01204277e-05 3.44068124e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381683e+00                   4
RALD3G                  C   3H   5O   1     G    300.00   3500.00 1160.00      1
-2.96412172e+00 3.83579385e-02-2.08581719e-05 5.12593560e-09-4.77571609e-13    2
 1.72028134e+03 4.58634919e+01 6.34826535e+00 6.24625900e-03 2.06655517e-05    3
-1.87382733e-08 4.66557687e-12-4.40192456e+02-4.45537170e-01                   4
RALDEST                 C   6H   9O   3     G    300.00   3500.00 1800.00      1
 1.17688624e+01 4.16586310e-02-2.02330626e-05 4.68126751e-09-4.21941087e-13    2
-4.91007178e+04-2.27507735e+01 5.76645054e+00 5.49973240e-02-3.13486401e-05    3
 8.79814806e-09-9.93730052e-13-4.69398496e+04 9.73553160e+00                   4
RBIPHENYL               C  12H   9          G    300.00   3500.00 1450.00      1
 2.67692078e+01 2.81611415e-02-6.05667723e-06-3.69378426e-10 1.67249382e-13    2
 3.92769947e+04-1.21306413e+02-1.05625108e+01 1.31145193e-01-1.12591903e-04    3
 4.86123345e-08-8.27787353e-12 5.01031931e+04 7.26686556e+01                   4
RBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1670.00      1
 1.45390319e+01 2.69797332e-02-1.09312485e-05 2.12602294e-09-1.64284673e-13    2
-3.56893368e+04-4.22613629e+01 3.26237571e+00 5.39896881e-02-3.51916871e-05    3
 1.18108288e-08-1.61410590e-12-3.19229337e+04 1.79249204e+01                   4
RC9H11                  C   9H  11          G    300.00   3500.00 1800.00      1
 1.94777671e+01 3.52558917e-02-1.42493230e-05 2.76058348e-09-2.13045169e-13    2
 6.10938819e+03-7.94713741e+01-1.83523003e+00 8.26181075e-02-5.37178363e-05    3
 1.73785513e-08-2.24331848e-12 1.37820672e+04 3.58790126e+01                   4
RCRESOLC                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541709e+01 2.50657189e-02-5.32353914e-06-2.12687585e-10 1.25840459e-13    2
-3.38086418e+03-4.22339552e+01-6.42956805e+00 9.31830717e-02-9.41722601e-05    3
 5.12938173e-08-1.10712258e-11 1.12339577e+03 5.49833259e+01                   4
RCRESOLO                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824813e+01 2.40796407e-02-4.51347946e-06-4.25076334e-10 1.44988488e-13    2
-3.97704754e+03-4.00543783e+01-6.60757189e+00 9.15233042e-02-9.24834752e-05    3
 5.05720227e-08-1.09413374e-11 4.82664709e+02 5.62014116e+01                   4
RDECALIN                C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278088e+00 9.04971362e+01                   4
RDECOO                  C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
RDIPE                   C   6H  13O   1     G    300.00   3500.00 1800.00      1
 1.69549494e+01 3.45118423e-02-1.31342732e-05 2.36150213e-09-1.67133125e-13    2
-2.78147477e+04-5.54607975e+01 6.91787207e-01 7.06522027e-02-4.32512401e-05    3
 1.35159343e-08-1.71635982e-12-2.19600093e+04 3.25588287e+01                   4
RMBOOX                  C   5H   9O   4     G    300.00   3500.00 1350.00      1
 2.46557066e+01 1.60203243e-02-2.33018024e-06-2.09432791e-10 5.96256606e-14    2
-5.87318865e+04-9.28197844e+01-3.02577545e+00 9.80395304e-02-9.34626315e-05    3
 4.47942468e-08-8.27438909e-12-5.12578864e+04 4.90347050e+01                   4
RMBX                    C   5H   9O   2     G    300.00   3500.00 1800.00      1
 1.54924702e+01 2.80794103e-02-1.20573254e-05 2.49322401e-09-2.04812728e-13    2
-3.97201864e+04-5.41810445e+01 2.13573311e+00 5.77610483e-02-3.67920237e-05    3
 1.16542234e-08-1.47717375e-12-3.49117610e+04 1.81084031e+01                   4
RMCROTA                 C   5H   7O   2     G    300.00   3500.00 1430.00      1
 1.57189282e+01 1.69463336e-02-4.46708252e-06 5.66631307e-10-2.76621493e-14    2
-3.23219582e+04-4.94508733e+01 1.47581476e-01 6.05025483e-02-5.01554196e-05    3
 2.18665554e-08-3.75142509e-12-2.78685530e+04 3.12413465e+01                   4
RMCYC6                  C   7H  13          G    300.00   3500.00 1800.00      1
 1.73339062e+01 3.85260822e-02-1.58310821e-05 3.15191459e-09-2.53163787e-13    2
-5.89957980e+03-7.33836419e+01-9.95790329e+00 9.91745477e-02-6.63714701e-05    3
 2.18705768e-08-2.85297798e-12 3.92547162e+03 7.43253244e+01                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.27624311e+01 3.77290665e-02-1.50512076e-05 2.88934934e-09-2.22140396e-13    2
-2.53740824e+04-9.90983226e+01-6.71698823e+00 1.03238887e-01-6.96427248e-05    3
 2.31084298e-08-3.03034602e-12-1.47614915e+04 6.04504445e+01                   4
RMDOOX                  C  11H  21O   4     G    300.00   3500.00 1800.00      1
 3.96894034e+01 5.38225057e-02-2.02775001e-05 3.64793874e-09-2.61216335e-13    2
-8.38472341e+04-1.67546736e+02 4.70466765e+00 1.31566363e-01-8.50640479e-05    3
 2.76429564e-08-3.59385768e-12-7.12527292e+04 2.17979520e+01                   4
RMDX                    C  11H  21O   2     G    300.00   3500.00 1800.00      1
 2.51620868e+01 7.14154614e-02-3.28250989e-05 7.27501997e-09-6.35222696e-13    2
-5.95987259e+04-9.23572595e+01 1.85440015e+00 1.23210321e-01-7.59874815e-05    3
 2.32610876e-08-2.85550987e-12-5.12079587e+04 3.37888029e+01                   4
RME7                    C   8H  15O   2     G    300.00   3500.00 1800.00      1
 2.40410392e+01 4.26053894e-02-1.71372001e-05 3.34440554e-09-2.61909734e-13    2
-4.89929735e+04-9.20931877e+01 2.93892065e+00 8.94989861e-02-5.62151974e-05    3
 1.78177379e-08-2.27209478e-12-4.13962109e+04 2.21158799e+01                   4
RMEOLEA                 C  19H  35O   2     G    300.00   3500.00 1800.00      1
 5.65772245e+01 8.98805970e-02-3.42288160e-05 6.24735813e-09-4.55216117e-13    2
-8.06885447e+04-2.49965378e+02-1.57106282e-01 2.15956888e-01-1.39292391e-04    3
 4.51597935e-08-5.85972103e-12-6.02641856e+04 5.70926555e+01                   4
RMEOLEOOX               C  19H  35O   4     G    300.00   3500.00 1800.00      1
 5.68288430e+01 9.87024571e-02-3.87236246e-05 7.19531442e-09-5.31279781e-13    2
-1.23280985e+05-2.44956753e+02 2.29713937e+00 2.19884021e-01-1.39708261e-04    3
 4.45970316e-08-5.72596272e-12-1.03649572e+05 5.01802030e+01                   4
RMEOLES                 C  19H  35O   2     G    300.00   3500.00 1800.00      1
 5.65772245e+01 8.98805970e-02-3.42288160e-05 6.24735813e-09-4.55216117e-13    2
-8.06885447e+04-2.49965378e+02-1.57106282e-01 2.15956888e-01-1.39292391e-04    3
 4.51597935e-08-5.85972103e-12-6.02641856e+04 5.70926555e+01                   4
RMLIN1A                 C  19H  31O   2     G    300.00   3500.00 1800.00      1
 5.95150691e+01 7.42461115e-02-2.53824843e-05 3.82833735e-09-2.08614643e-13    2
-4.82863749e+04-2.69048825e+02-9.12524230e-01 2.08529652e-01-1.37285435e-04    3
 4.52738746e-08-5.96493926e-12-2.65324413e+04 5.79979154e+01                   4
RMLIN1OOX               C  19H  31O   4     G    300.00   3500.00 1650.00      1
 5.48798863e+01 9.05843840e-02-3.54321193e-05 6.50176029e-09-4.69049023e-13    2
-7.13229393e+04-2.34809039e+02-1.47497564e+00 2.27202231e-01-1.59630162e-04    3
 5.66827877e-08-8.07223499e-12-5.27258349e+04 6.52917158e+01                   4
RMLIN1X                 C  19H  31O   2     G    300.00   3500.00 1800.00      1
 5.95150691e+01 7.42461115e-02-2.53824843e-05 3.82833735e-09-2.08614643e-13    2
-4.82863749e+04-2.69048825e+02-9.12524230e-01 2.08529652e-01-1.37285435e-04    3
 4.52738746e-08-5.96493926e-12-2.65324413e+04 5.79979154e+01                   4
RMLINA                  C  19H  33O   2     G    300.00   3500.00 1800.00      1
 5.71954712e+01 8.40022248e-02-3.15645422e-05 5.64019755e-09-4.00096883e-13    2
-6.69574846e+04-2.54485602e+02-1.30856133e+00 2.14011186e-01-1.39905343e-04    3
 4.57664202e-08-5.97318336e-12-4.58960329e+04 6.21504271e+01                   4
RMLINOOX                C  19H  33O   4     G    300.00   3500.00 1780.00      1
 6.32132444e+01 8.05239356e-02-2.78197745e-05 4.27200724e-09-2.39927804e-13    2
-8.77238917e+04-2.82700411e+02 1.99661323e+00 2.18089399e-01-1.43745727e-04    3
 4.76899669e-08-6.33795584e-12-6.59307710e+04 4.79327752e+01                   4
RMLINX                  C  19H  33O   2     G    300.00   3500.00 1800.00      1
 5.71954712e+01 8.40022248e-02-3.15645422e-05 5.64019755e-09-4.00096883e-13    2
-6.69574846e+04-2.54485602e+02-1.30856133e+00 2.14011186e-01-1.39905343e-04    3
 4.57664202e-08-5.97318336e-12-4.58960329e+04 6.21504271e+01                   4
RMP3                    C   4H   7O   2     G    300.00   3500.00 1800.00      1
 9.46731146e+00 2.78903391e-02-1.31079861e-05 2.94998316e-09-2.60075548e-13    2
-3.18264551e+04-1.93081295e+01 3.67472870e+00 4.07627453e-02-2.38349912e-05    3
 6.92294802e-09-8.11876222e-13-2.97411253e+04 1.20425368e+01                   4
RMPAOOX                 C  17H  33O   4     G    300.00   3500.00 1800.00      1
 3.96894034e+01 5.38225057e-02-2.02775001e-05 3.64793874e-09-2.61216335e-13    2
-8.38472341e+04-1.67546736e+02 4.70466765e+00 1.31566363e-01-8.50640479e-05    3
 2.76429564e-08-3.59385768e-12-7.12527292e+04 2.17979520e+01                   4
RMPAX                   C  17H  33O   2     G    300.00   3500.00 1570.00      1
 4.65991944e+01 8.79958559e-02-3.11818152e-05 4.72867036e-09-2.34133930e-13    2
-8.86750528e+04-2.03460488e+02-5.53001427e+00 2.20809126e-01-1.58073475e-04    3
 5.86104792e-08-8.81403979e-12-7.23064813e+04 7.15470253e+01                   4
RMSTEAOOX               C  19H  37O   4     G    300.00   3500.00 1250.00      1
-1.20700825e+02 5.67736647e-01-4.52750605e-04 1.47317719e-07-1.67528750e-11    2
 1.02039730e+04 6.60024010e+02 1.91170969e+01 1.20319297e-01 8.41502162e-05    3
-1.39029386e-07 4.05165459e-11-2.47505076e+04-4.57161098e+01                   4
RMTBE                   C   5H  11O   1     G    300.00   3500.00 1370.00      1
 1.09269229e+01 3.74766266e-02-1.73062474e-05 3.86241414e-09-3.39119741e-13    2
-1.88007827e+04-2.53563680e+01-1.81069448e-01 6.99087211e-02-5.28158399e-05    3
 2.11420212e-08-3.49233271e-12-1.57571928e+04 3.17301895e+01                   4
RODECA                  C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278088e+00 9.04971362e+01                   4
RSTEAX                  C  19H  37O   2     G    300.00   3500.00 1590.00      1
 5.46335802e+01 9.34230719e-02-3.19964312e-05 4.67181818e-09-2.16706943e-13    2
-9.74617261e+04-2.43777088e+02-6.34709308e+00 2.46833571e-01-1.76723317e-04    3
 6.53539506e-08-9.75792273e-12-7.80698720e+04 7.86982236e+01                   4
RTC4H8OH                C   4H   9O   1     G    300.00   3500.00 1380.00      1
 8.66823484e+00 3.01271731e-02-1.35256253e-05 2.94117291e-09-2.52822189e-13    2
-1.73478965e+04-1.68023720e+01 1.39901320e-03 5.52484364e-02-4.08313463e-05    3
 1.61323424e-08-2.64252681e-12-1.49558499e+04 2.78015457e+01                   4
RTC4H9O                 C   4H   9O   1     G    300.00   3500.00 1610.00      1
 1.16852527e+01 2.57155374e-02-1.07539562e-05 2.15924613e-09-1.71897014e-13    2
-1.72607591e+04-3.73085633e+01-2.94435988e-01 5.54787390e-02-3.84836472e-05    3
 1.36415198e-08-1.95485877e-12-1.34032994e+04 2.61916467e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92428061e+01 2.67835937e-02-9.17249482e-06 1.42952536e-09-8.46466186e-14    2
 3.95646504e+03-1.44540610e+02-1.09331575e+01 1.16063513e-01-8.35724273e-05    3
 2.89850559e-08-3.91180364e-12 1.84198119e+04 7.29000859e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619031e+01-7.89283132e-03 1.09697206e-05-3.89489830e-09 4.38586293e-13    2
-1.76924159e+04-2.71823424e+02-1.36343924e+01 1.41210048e-01-1.13282678e-04    3
 4.21245088e-08-5.95299802e-12 6.46225047e+03 9.13157248e+01                   4
RUME10                  C  11H  19O   2     G    300.00   3500.00 1450.00      1
 2.35916369e+01 6.52041736e-02-2.68467537e-05 5.44034955e-09-4.42864735e-13    2
-3.58672705e+04-8.27430018e+01 1.64400814e+00 1.25749356e-01-8.94797013e-05    3
 3.42371070e-08-5.40782293e-12-2.95024582e+04 3.12965588e+01                   4
RUME16                  C  17H  31O   2     G    300.00   3500.00 1790.00      1
 5.62816009e+01 7.14355580e-02-2.43272135e-05 3.65699376e-09-1.98260551e-13    2
-7.53409955e+04-2.53924384e+02 9.94524607e-01 1.94982097e-01-1.27857833e-04    3
 4.22158836e-08-5.58358037e-12-5.55482222e+04 4.49927995e+01                   4
RUME7                   C   8H  13O   2     G    300.00   3500.00 1800.00      1
 1.85903431e+01 4.63199659e-02-2.12076343e-05 4.67919597e-09-4.06994657e-13    2
-3.29183962e+04-6.07637830e+01 2.66158720e+00 8.17172013e-02-5.07053305e-05    3
 1.56042686e-08-1.92436586e-12-2.71840440e+04 2.54459670e+01                   4
RXYLENE                 C   8H   9          G    300.00   3500.00 1380.00      1
 9.50606195e+00 4.15939315e-02-1.79471777e-05 3.41861978e-09-2.36020443e-13    2
 1.46969060e+04-2.59567399e+01-2.80920460e+00 7.72903563e-02-5.67476394e-05    3
 2.21628042e-08-3.63170602e-12 1.80959195e+04 3.74238465e+01                   4
SC4H7                   C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017753e+00 1.98466503e-02-6.37614062e-06 5.28652771e-10 3.81103730e-14    2
 1.19533850e+04-1.83767118e+01-1.12550124e+00 4.64823652e-02-3.45124591e-05    3
 1.37381920e-08-2.28751273e-12 1.46387978e+04 3.05571711e+01                   4
TAME                    C   6H  14O   1     G    300.00   3500.00 1320.00      1
 1.13309761e+01 4.74280944e-02-1.96957502e-05 3.66860750e-09-2.50688228e-13    2
-4.42745214e+04-3.17952394e+01-2.12836721e+00 8.82139832e-02-6.60433511e-05    3
 2.70764868e-08-4.68399869e-12-4.07212548e+04 3.68750527e+01                   4
TC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1440.00      1
 9.08150387e+00 3.22201837e-02-1.41979352e-05 3.03249263e-09-2.56658356e-13    2
-4.23917231e+04-2.36263218e+01-6.99999563e-01 5.93910266e-02-4.25008966e-05    3
 1.61357155e-08-2.53152343e-12-3.95746501e+04 2.71305359e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250678e+01 3.45031690e-02-1.26565536e-05 2.20632462e-09-1.51941206e-13    2
-9.85314330e+03-1.11161769e+02-1.00807336e+01 1.17183900e-01-8.78208542e-05    3
 3.25757390e-08-4.75336763e-12 1.40177116e+03 7.04583499e+01                   4
TMBENZ                  C   9H  12          G    300.00   3500.00 1800.00      1
 1.47576861e+01 4.50315825e-02-1.97554195e-05 4.21197817e-09-3.57314917e-13    2
-1.09025839e+04-5.35378398e+01-2.75522789e+00 8.39491691e-02-5.21867417e-05    3
 1.62235790e-08-2.02559281e-12-4.59793488e+03 4.12457040e+01                   4
U2ME10                  C  11H  18O   2     G    300.00   3500.00 1440.00      1
 2.36788649e+01 6.40632046e-02-2.76021386e-05 5.83270375e-09-4.91952687e-13    2
-5.39118596e+04-8.57548642e+01 3.22839337e-01 1.28941053e-01-9.51832310e-05    3
 3.71202465e-08-5.92381775e-12-4.71853243e+04 3.54410717e+01                   4
U2ME12                  C  13H  22O   2     G    300.00   3500.00 1610.00      1
 3.12799449e+01 7.15415882e-02-3.01181538e-05 6.08643201e-09-4.87334868e-13    2
-6.28268100e+04-1.24478592e+02 1.12650720e+00 1.46456961e-01-9.99150853e-05    3
 3.49878529e-08-4.97513315e-12-5.31174030e+04 3.53544123e+01                   4
UME10                   C  11H  20O   2     G    300.00   3500.00 1800.00      1
 3.48566736e+01 5.08631615e-02-1.90027410e-05 3.39432106e-09-2.41664061e-13    2
-7.27334602e+04-1.48477392e+02 1.08700033e+00 1.25906880e-01-8.15391729e-05    3
 2.65559625e-08-3.45855871e-12-6.05763778e+04 3.42911241e+01                   4
UME16                   C  17H  32O   2     G    300.00   3500.00 1580.00      1
 4.52339702e+01 8.65152352e-02-3.05153342e-05 4.60674378e-09-2.26752205e-13    2
-9.22046847e+04-1.94026893e+02-6.34895832e+00 2.17104928e-01-1.54492890e-04    3
 5.69179489e-08-8.50384163e-12-7.59044793e+04 7.84262324e+01                   4
UME7                    C   8H  14O   2     G    300.00   3500.00 1800.00      1
 2.58473842e+01 3.62113327e-02-1.33124030e-05 2.32937526e-09-1.61944568e-13    2
-5.91274188e+04-1.03960065e+02 2.21977808e+00 8.87171241e-02-5.70672292e-05    3
 1.85348664e-08-2.41270723e-12-5.06214805e+04 2.39174684e+01                   4
XYLENE                  C   8H  10          G    300.00   3500.00 1640.00      1
 1.72256243e+01 2.83565600e-02-6.90689954e-06-3.57091403e-10 2.09419626e-13    2
-6.87239337e+03-6.97341599e+01-5.12303971e+00 8.28654966e-02-5.67626342e-05    3
 1.99094674e-08-2.87999483e-12 4.57968429e+02 4.91410252e+01                   4
ZBU1OOX                 C   4H   9O   5     G    300.00   3500.00 1410.00      1
 1.71509971e+01 3.21642995e-02-1.45265250e-05 3.16055984e-09-2.71089893e-13    2
-4.87167967e+04-4.94521678e+01 4.90929016e+00 6.68925461e-02-5.14714682e-05    3
 2.06286181e-08-3.36826334e-12-4.52646353e+04 1.38131161e+01                   4
ZDECA                   C  10H  17O   4     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
ZMBOOX                  C   5H   9O   6     G    300.00   3500.00 1310.00      1
 2.94016942e+01 1.57346453e-02-2.10565670e-06-2.30310175e-10 5.80528651e-14    2
-7.03637113e+04-1.09596841e+02-1.66570869e+00 1.10596944e-01-1.10726610e-04    3
 5.50475284e-08-1.04911530e-11-6.22240518e+04 4.86744607e+01                   4
ZMDOOH                  C  11H  21O   6     G    300.00   3500.00 1780.00      1
 4.89601122e+01 4.69646617e-02-1.61477773e-05 2.58757356e-09-1.58080023e-13    2
-9.96313675e+04-2.11226530e+02 6.91495056e+00 1.41448171e-01-9.57687121e-05    3
 3.24081484e-08-4.34636300e-12-8.46632899e+04 1.58608722e+01                   4
ZMEOLEOOX               C  19H  35O   6     G    300.00   3500.00 1540.00      1
 5.74950108e+01 9.92606422e-02-3.35004082e-05 5.08063679e-09-2.82240300e-13    2
-1.09648465e+05-2.38315353e+02 2.38451828e+00 2.42404779e-01-1.72926515e-04    3
 6.54382588e-08-1.00805556e-11-9.26744334e+04 5.13566583e+01                   4
ZMLIN1OOX               C  19H  31O   6     G    300.00   3500.00 1690.00      1
 6.61920071e+01 8.18444133e-02-3.03706056e-05 5.17171152e-09-3.39000627e-13    2
-8.83104294e+04-2.93138255e+02 7.95447186e-01 2.36629171e-01-1.67753526e-04    3
 5.93661575e-08-8.35593051e-12-6.62063921e+04 5.66777851e+01                   4
ZMLINOOX                C  19H  33O   6     G    300.00   3500.00 1530.00      1
 6.14087077e+01 8.58331824e-02-2.98017595e-05 4.63939709e-09-2.65661024e-13    2
-9.65914210e+04-2.81173958e+02 1.31186651e+00 2.42949107e-01-1.83836980e-04    3
 7.17571402e-08-1.12326125e-11-7.82017876e+04 3.43158089e+01                   4
ZMPAOOH                 C  17H  33O   6     G    300.00   3500.00 1780.00      1
 4.89601122e+01 4.69646617e-02-1.61477773e-05 2.58757356e-09-1.58080023e-13    2
-9.96313675e+04-2.11226530e+02 6.91495056e+00 1.41448171e-01-9.57687121e-05    3
 3.24081484e-08-4.34636300e-12-8.46632899e+04 1.58608722e+01                   4
ZMSTEAOOH               C  19H  37O   6     G    300.00   3500.00 1250.00      1
-6.22995292e+01 3.41575945e-01-2.69706994e-04 8.71969173e-08-9.87435445e-12    2
 1.57160052e+04 3.57020399e+02 1.61954271e+01 9.03920846e-02 3.17136382e-05    3
-7.35607531e-08 2.22771796e-11-3.90773390e+03-3.91880337e+01                   4
END
